//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Top-level Verilog module for FPGA
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Mon Dec  9 17:13:32 2024
//-------------------------------------------
//----- Time scale -----
`timescale 1ns / 1ps

//----- Default net type -----
`default_nettype wire

// ----- Verilog module for fpga_top -----
module fpga_top(clk,
                reset,
                isol_n,
                pReset,
                prog_clk,
                Test_en,
                gfpga_pad_io_soc_in,
                gfpga_pad_io_soc_out,
                gfpga_pad_io_soc_dir,
                ccff_head,
                ccff_tail);
//----- GLOBAL PORTS -----
input [0:0] clk;
//----- GLOBAL PORTS -----
input [0:0] reset;
//----- GLOBAL PORTS -----
input [0:0] isol_n;
//----- GLOBAL PORTS -----
input [0:0] pReset;
//----- GLOBAL PORTS -----
input [0:0] prog_clk;
//----- GLOBAL PORTS -----
input [0:0] Test_en;
//----- GPIN PORTS -----
input [0:127] gfpga_pad_io_soc_in;
//----- GPOUT PORTS -----
output [0:127] gfpga_pad_io_soc_out;
//----- GPOUT PORTS -----
output [0:127] gfpga_pad_io_soc_dir;
//----- INPUT PORTS -----
input [0:0] ccff_head;
//----- OUTPUT PORTS -----
output [0:0] ccff_tail;

//----- BEGIN Registered ports -----
//----- END Registered ports -----


wire [0:29] cbx_1__0__0_chanx_left_out;
wire [0:29] cbx_1__0__0_chanx_right_out;
wire [0:29] cbx_1__0__1_chanx_left_out;
wire [0:29] cbx_1__0__1_chanx_right_out;
wire [0:29] cbx_1__0__2_chanx_left_out;
wire [0:29] cbx_1__0__2_chanx_right_out;
wire [0:29] cbx_1__0__3_chanx_left_out;
wire [0:29] cbx_1__0__3_chanx_right_out;
wire [0:29] cbx_1__0__4_chanx_left_out;
wire [0:29] cbx_1__0__4_chanx_right_out;
wire [0:29] cbx_1__0__5_chanx_left_out;
wire [0:29] cbx_1__0__5_chanx_right_out;
wire [0:29] cbx_1__0__6_chanx_left_out;
wire [0:29] cbx_1__0__6_chanx_right_out;
wire [0:29] cbx_1__0__7_chanx_left_out;
wire [0:29] cbx_1__0__7_chanx_right_out;
wire [0:29] cbx_1__1__0_chanx_left_out;
wire [0:29] cbx_1__1__0_chanx_right_out;
wire [0:29] cbx_1__1__10_chanx_left_out;
wire [0:29] cbx_1__1__10_chanx_right_out;
wire [0:29] cbx_1__1__11_chanx_left_out;
wire [0:29] cbx_1__1__11_chanx_right_out;
wire [0:29] cbx_1__1__12_chanx_left_out;
wire [0:29] cbx_1__1__12_chanx_right_out;
wire [0:29] cbx_1__1__13_chanx_left_out;
wire [0:29] cbx_1__1__13_chanx_right_out;
wire [0:29] cbx_1__1__14_chanx_left_out;
wire [0:29] cbx_1__1__14_chanx_right_out;
wire [0:29] cbx_1__1__15_chanx_left_out;
wire [0:29] cbx_1__1__15_chanx_right_out;
wire [0:29] cbx_1__1__16_chanx_left_out;
wire [0:29] cbx_1__1__16_chanx_right_out;
wire [0:29] cbx_1__1__17_chanx_left_out;
wire [0:29] cbx_1__1__17_chanx_right_out;
wire [0:29] cbx_1__1__18_chanx_left_out;
wire [0:29] cbx_1__1__18_chanx_right_out;
wire [0:29] cbx_1__1__19_chanx_left_out;
wire [0:29] cbx_1__1__19_chanx_right_out;
wire [0:29] cbx_1__1__1_chanx_left_out;
wire [0:29] cbx_1__1__1_chanx_right_out;
wire [0:29] cbx_1__1__20_chanx_left_out;
wire [0:29] cbx_1__1__20_chanx_right_out;
wire [0:29] cbx_1__1__21_chanx_left_out;
wire [0:29] cbx_1__1__21_chanx_right_out;
wire [0:29] cbx_1__1__22_chanx_left_out;
wire [0:29] cbx_1__1__22_chanx_right_out;
wire [0:29] cbx_1__1__23_chanx_left_out;
wire [0:29] cbx_1__1__23_chanx_right_out;
wire [0:29] cbx_1__1__24_chanx_left_out;
wire [0:29] cbx_1__1__24_chanx_right_out;
wire [0:29] cbx_1__1__25_chanx_left_out;
wire [0:29] cbx_1__1__25_chanx_right_out;
wire [0:29] cbx_1__1__26_chanx_left_out;
wire [0:29] cbx_1__1__26_chanx_right_out;
wire [0:29] cbx_1__1__27_chanx_left_out;
wire [0:29] cbx_1__1__27_chanx_right_out;
wire [0:29] cbx_1__1__28_chanx_left_out;
wire [0:29] cbx_1__1__28_chanx_right_out;
wire [0:29] cbx_1__1__29_chanx_left_out;
wire [0:29] cbx_1__1__29_chanx_right_out;
wire [0:29] cbx_1__1__2_chanx_left_out;
wire [0:29] cbx_1__1__2_chanx_right_out;
wire [0:29] cbx_1__1__30_chanx_left_out;
wire [0:29] cbx_1__1__30_chanx_right_out;
wire [0:29] cbx_1__1__31_chanx_left_out;
wire [0:29] cbx_1__1__31_chanx_right_out;
wire [0:29] cbx_1__1__32_chanx_left_out;
wire [0:29] cbx_1__1__32_chanx_right_out;
wire [0:29] cbx_1__1__33_chanx_left_out;
wire [0:29] cbx_1__1__33_chanx_right_out;
wire [0:29] cbx_1__1__34_chanx_left_out;
wire [0:29] cbx_1__1__34_chanx_right_out;
wire [0:29] cbx_1__1__35_chanx_left_out;
wire [0:29] cbx_1__1__35_chanx_right_out;
wire [0:29] cbx_1__1__36_chanx_left_out;
wire [0:29] cbx_1__1__36_chanx_right_out;
wire [0:29] cbx_1__1__37_chanx_left_out;
wire [0:29] cbx_1__1__37_chanx_right_out;
wire [0:29] cbx_1__1__38_chanx_left_out;
wire [0:29] cbx_1__1__38_chanx_right_out;
wire [0:29] cbx_1__1__39_chanx_left_out;
wire [0:29] cbx_1__1__39_chanx_right_out;
wire [0:29] cbx_1__1__3_chanx_left_out;
wire [0:29] cbx_1__1__3_chanx_right_out;
wire [0:29] cbx_1__1__40_chanx_left_out;
wire [0:29] cbx_1__1__40_chanx_right_out;
wire [0:29] cbx_1__1__41_chanx_left_out;
wire [0:29] cbx_1__1__41_chanx_right_out;
wire [0:29] cbx_1__1__42_chanx_left_out;
wire [0:29] cbx_1__1__42_chanx_right_out;
wire [0:29] cbx_1__1__43_chanx_left_out;
wire [0:29] cbx_1__1__43_chanx_right_out;
wire [0:29] cbx_1__1__44_chanx_left_out;
wire [0:29] cbx_1__1__44_chanx_right_out;
wire [0:29] cbx_1__1__45_chanx_left_out;
wire [0:29] cbx_1__1__45_chanx_right_out;
wire [0:29] cbx_1__1__46_chanx_left_out;
wire [0:29] cbx_1__1__46_chanx_right_out;
wire [0:29] cbx_1__1__47_chanx_left_out;
wire [0:29] cbx_1__1__47_chanx_right_out;
wire [0:29] cbx_1__1__48_chanx_left_out;
wire [0:29] cbx_1__1__48_chanx_right_out;
wire [0:29] cbx_1__1__49_chanx_left_out;
wire [0:29] cbx_1__1__49_chanx_right_out;
wire [0:29] cbx_1__1__4_chanx_left_out;
wire [0:29] cbx_1__1__4_chanx_right_out;
wire [0:29] cbx_1__1__50_chanx_left_out;
wire [0:29] cbx_1__1__50_chanx_right_out;
wire [0:29] cbx_1__1__51_chanx_left_out;
wire [0:29] cbx_1__1__51_chanx_right_out;
wire [0:29] cbx_1__1__52_chanx_left_out;
wire [0:29] cbx_1__1__52_chanx_right_out;
wire [0:29] cbx_1__1__53_chanx_left_out;
wire [0:29] cbx_1__1__53_chanx_right_out;
wire [0:29] cbx_1__1__54_chanx_left_out;
wire [0:29] cbx_1__1__54_chanx_right_out;
wire [0:29] cbx_1__1__55_chanx_left_out;
wire [0:29] cbx_1__1__55_chanx_right_out;
wire [0:29] cbx_1__1__5_chanx_left_out;
wire [0:29] cbx_1__1__5_chanx_right_out;
wire [0:29] cbx_1__1__6_chanx_left_out;
wire [0:29] cbx_1__1__6_chanx_right_out;
wire [0:29] cbx_1__1__7_chanx_left_out;
wire [0:29] cbx_1__1__7_chanx_right_out;
wire [0:29] cbx_1__1__8_chanx_left_out;
wire [0:29] cbx_1__1__8_chanx_right_out;
wire [0:29] cbx_1__1__9_chanx_left_out;
wire [0:29] cbx_1__1__9_chanx_right_out;
wire [0:29] cbx_1__8__0_chanx_left_out;
wire [0:29] cbx_1__8__0_chanx_right_out;
wire [0:29] cbx_1__8__1_chanx_left_out;
wire [0:29] cbx_1__8__1_chanx_right_out;
wire [0:29] cbx_1__8__2_chanx_left_out;
wire [0:29] cbx_1__8__2_chanx_right_out;
wire [0:29] cbx_1__8__3_chanx_left_out;
wire [0:29] cbx_1__8__3_chanx_right_out;
wire [0:29] cbx_1__8__4_chanx_left_out;
wire [0:29] cbx_1__8__4_chanx_right_out;
wire [0:29] cbx_1__8__5_chanx_left_out;
wire [0:29] cbx_1__8__5_chanx_right_out;
wire [0:29] cbx_1__8__6_chanx_left_out;
wire [0:29] cbx_1__8__6_chanx_right_out;
wire [0:29] cbx_1__8__7_chanx_left_out;
wire [0:29] cbx_1__8__7_chanx_right_out;
wire [0:29] cby_0__1__0_chany_bottom_out;
wire [0:29] cby_0__1__0_chany_top_out;
wire [0:29] cby_0__1__1_chany_bottom_out;
wire [0:29] cby_0__1__1_chany_top_out;
wire [0:29] cby_0__1__2_chany_bottom_out;
wire [0:29] cby_0__1__2_chany_top_out;
wire [0:29] cby_0__1__3_chany_bottom_out;
wire [0:29] cby_0__1__3_chany_top_out;
wire [0:29] cby_0__1__4_chany_bottom_out;
wire [0:29] cby_0__1__4_chany_top_out;
wire [0:29] cby_0__1__5_chany_bottom_out;
wire [0:29] cby_0__1__5_chany_top_out;
wire [0:29] cby_0__1__6_chany_bottom_out;
wire [0:29] cby_0__1__6_chany_top_out;
wire [0:29] cby_0__1__7_chany_bottom_out;
wire [0:29] cby_0__1__7_chany_top_out;
wire [0:29] cby_1__1__0_chany_bottom_out;
wire [0:29] cby_1__1__0_chany_top_out;
wire [0:29] cby_1__1__10_chany_bottom_out;
wire [0:29] cby_1__1__10_chany_top_out;
wire [0:29] cby_1__1__11_chany_bottom_out;
wire [0:29] cby_1__1__11_chany_top_out;
wire [0:29] cby_1__1__12_chany_bottom_out;
wire [0:29] cby_1__1__12_chany_top_out;
wire [0:29] cby_1__1__13_chany_bottom_out;
wire [0:29] cby_1__1__13_chany_top_out;
wire [0:29] cby_1__1__14_chany_bottom_out;
wire [0:29] cby_1__1__14_chany_top_out;
wire [0:29] cby_1__1__15_chany_bottom_out;
wire [0:29] cby_1__1__15_chany_top_out;
wire [0:29] cby_1__1__16_chany_bottom_out;
wire [0:29] cby_1__1__16_chany_top_out;
wire [0:29] cby_1__1__17_chany_bottom_out;
wire [0:29] cby_1__1__17_chany_top_out;
wire [0:29] cby_1__1__18_chany_bottom_out;
wire [0:29] cby_1__1__18_chany_top_out;
wire [0:29] cby_1__1__19_chany_bottom_out;
wire [0:29] cby_1__1__19_chany_top_out;
wire [0:29] cby_1__1__1_chany_bottom_out;
wire [0:29] cby_1__1__1_chany_top_out;
wire [0:29] cby_1__1__20_chany_bottom_out;
wire [0:29] cby_1__1__20_chany_top_out;
wire [0:29] cby_1__1__21_chany_bottom_out;
wire [0:29] cby_1__1__21_chany_top_out;
wire [0:29] cby_1__1__22_chany_bottom_out;
wire [0:29] cby_1__1__22_chany_top_out;
wire [0:29] cby_1__1__23_chany_bottom_out;
wire [0:29] cby_1__1__23_chany_top_out;
wire [0:29] cby_1__1__24_chany_bottom_out;
wire [0:29] cby_1__1__24_chany_top_out;
wire [0:29] cby_1__1__25_chany_bottom_out;
wire [0:29] cby_1__1__25_chany_top_out;
wire [0:29] cby_1__1__26_chany_bottom_out;
wire [0:29] cby_1__1__26_chany_top_out;
wire [0:29] cby_1__1__27_chany_bottom_out;
wire [0:29] cby_1__1__27_chany_top_out;
wire [0:29] cby_1__1__28_chany_bottom_out;
wire [0:29] cby_1__1__28_chany_top_out;
wire [0:29] cby_1__1__29_chany_bottom_out;
wire [0:29] cby_1__1__29_chany_top_out;
wire [0:29] cby_1__1__2_chany_bottom_out;
wire [0:29] cby_1__1__2_chany_top_out;
wire [0:29] cby_1__1__30_chany_bottom_out;
wire [0:29] cby_1__1__30_chany_top_out;
wire [0:29] cby_1__1__31_chany_bottom_out;
wire [0:29] cby_1__1__31_chany_top_out;
wire [0:29] cby_1__1__32_chany_bottom_out;
wire [0:29] cby_1__1__32_chany_top_out;
wire [0:29] cby_1__1__33_chany_bottom_out;
wire [0:29] cby_1__1__33_chany_top_out;
wire [0:29] cby_1__1__34_chany_bottom_out;
wire [0:29] cby_1__1__34_chany_top_out;
wire [0:29] cby_1__1__35_chany_bottom_out;
wire [0:29] cby_1__1__35_chany_top_out;
wire [0:29] cby_1__1__36_chany_bottom_out;
wire [0:29] cby_1__1__36_chany_top_out;
wire [0:29] cby_1__1__37_chany_bottom_out;
wire [0:29] cby_1__1__37_chany_top_out;
wire [0:29] cby_1__1__38_chany_bottom_out;
wire [0:29] cby_1__1__38_chany_top_out;
wire [0:29] cby_1__1__39_chany_bottom_out;
wire [0:29] cby_1__1__39_chany_top_out;
wire [0:29] cby_1__1__3_chany_bottom_out;
wire [0:29] cby_1__1__3_chany_top_out;
wire [0:29] cby_1__1__40_chany_bottom_out;
wire [0:29] cby_1__1__40_chany_top_out;
wire [0:29] cby_1__1__41_chany_bottom_out;
wire [0:29] cby_1__1__41_chany_top_out;
wire [0:29] cby_1__1__42_chany_bottom_out;
wire [0:29] cby_1__1__42_chany_top_out;
wire [0:29] cby_1__1__43_chany_bottom_out;
wire [0:29] cby_1__1__43_chany_top_out;
wire [0:29] cby_1__1__44_chany_bottom_out;
wire [0:29] cby_1__1__44_chany_top_out;
wire [0:29] cby_1__1__45_chany_bottom_out;
wire [0:29] cby_1__1__45_chany_top_out;
wire [0:29] cby_1__1__46_chany_bottom_out;
wire [0:29] cby_1__1__46_chany_top_out;
wire [0:29] cby_1__1__47_chany_bottom_out;
wire [0:29] cby_1__1__47_chany_top_out;
wire [0:29] cby_1__1__48_chany_bottom_out;
wire [0:29] cby_1__1__48_chany_top_out;
wire [0:29] cby_1__1__49_chany_bottom_out;
wire [0:29] cby_1__1__49_chany_top_out;
wire [0:29] cby_1__1__4_chany_bottom_out;
wire [0:29] cby_1__1__4_chany_top_out;
wire [0:29] cby_1__1__50_chany_bottom_out;
wire [0:29] cby_1__1__50_chany_top_out;
wire [0:29] cby_1__1__51_chany_bottom_out;
wire [0:29] cby_1__1__51_chany_top_out;
wire [0:29] cby_1__1__52_chany_bottom_out;
wire [0:29] cby_1__1__52_chany_top_out;
wire [0:29] cby_1__1__53_chany_bottom_out;
wire [0:29] cby_1__1__53_chany_top_out;
wire [0:29] cby_1__1__54_chany_bottom_out;
wire [0:29] cby_1__1__54_chany_top_out;
wire [0:29] cby_1__1__55_chany_bottom_out;
wire [0:29] cby_1__1__55_chany_top_out;
wire [0:29] cby_1__1__5_chany_bottom_out;
wire [0:29] cby_1__1__5_chany_top_out;
wire [0:29] cby_1__1__6_chany_bottom_out;
wire [0:29] cby_1__1__6_chany_top_out;
wire [0:29] cby_1__1__7_chany_bottom_out;
wire [0:29] cby_1__1__7_chany_top_out;
wire [0:29] cby_1__1__8_chany_bottom_out;
wire [0:29] cby_1__1__8_chany_top_out;
wire [0:29] cby_1__1__9_chany_bottom_out;
wire [0:29] cby_1__1__9_chany_top_out;
wire [0:29] cby_8__1__0_chany_bottom_out;
wire [0:29] cby_8__1__0_chany_top_out;
wire [0:29] cby_8__1__1_chany_bottom_out;
wire [0:29] cby_8__1__1_chany_top_out;
wire [0:29] cby_8__1__2_chany_bottom_out;
wire [0:29] cby_8__1__2_chany_top_out;
wire [0:29] cby_8__1__3_chany_bottom_out;
wire [0:29] cby_8__1__3_chany_top_out;
wire [0:29] cby_8__1__4_chany_bottom_out;
wire [0:29] cby_8__1__4_chany_top_out;
wire [0:29] cby_8__1__5_chany_bottom_out;
wire [0:29] cby_8__1__5_chany_top_out;
wire [0:29] cby_8__1__6_chany_bottom_out;
wire [0:29] cby_8__1__6_chany_top_out;
wire [0:29] cby_8__1__7_chany_bottom_out;
wire [0:29] cby_8__1__7_chany_top_out;
wire [0:29] sb_0__0__0_chanx_right_out;
wire [0:29] sb_0__0__0_chany_top_out;
wire [0:29] sb_0__1__0_chanx_right_out;
wire [0:29] sb_0__1__0_chany_bottom_out;
wire [0:29] sb_0__1__0_chany_top_out;
wire [0:29] sb_0__1__1_chanx_right_out;
wire [0:29] sb_0__1__1_chany_bottom_out;
wire [0:29] sb_0__1__1_chany_top_out;
wire [0:29] sb_0__1__2_chanx_right_out;
wire [0:29] sb_0__1__2_chany_bottom_out;
wire [0:29] sb_0__1__2_chany_top_out;
wire [0:29] sb_0__1__3_chanx_right_out;
wire [0:29] sb_0__1__3_chany_bottom_out;
wire [0:29] sb_0__1__3_chany_top_out;
wire [0:29] sb_0__1__4_chanx_right_out;
wire [0:29] sb_0__1__4_chany_bottom_out;
wire [0:29] sb_0__1__4_chany_top_out;
wire [0:29] sb_0__1__5_chanx_right_out;
wire [0:29] sb_0__1__5_chany_bottom_out;
wire [0:29] sb_0__1__5_chany_top_out;
wire [0:29] sb_0__1__6_chanx_right_out;
wire [0:29] sb_0__1__6_chany_bottom_out;
wire [0:29] sb_0__1__6_chany_top_out;
wire [0:29] sb_0__8__0_chanx_right_out;
wire [0:29] sb_0__8__0_chany_bottom_out;
wire [0:29] sb_1__0__0_chanx_left_out;
wire [0:29] sb_1__0__0_chanx_right_out;
wire [0:29] sb_1__0__0_chany_top_out;
wire [0:29] sb_1__0__1_chanx_left_out;
wire [0:29] sb_1__0__1_chanx_right_out;
wire [0:29] sb_1__0__1_chany_top_out;
wire [0:29] sb_1__0__2_chanx_left_out;
wire [0:29] sb_1__0__2_chanx_right_out;
wire [0:29] sb_1__0__2_chany_top_out;
wire [0:29] sb_1__0__3_chanx_left_out;
wire [0:29] sb_1__0__3_chanx_right_out;
wire [0:29] sb_1__0__3_chany_top_out;
wire [0:29] sb_1__0__4_chanx_left_out;
wire [0:29] sb_1__0__4_chanx_right_out;
wire [0:29] sb_1__0__4_chany_top_out;
wire [0:29] sb_1__0__5_chanx_left_out;
wire [0:29] sb_1__0__5_chanx_right_out;
wire [0:29] sb_1__0__5_chany_top_out;
wire [0:29] sb_1__0__6_chanx_left_out;
wire [0:29] sb_1__0__6_chanx_right_out;
wire [0:29] sb_1__0__6_chany_top_out;
wire [0:29] sb_1__1__0_chanx_left_out;
wire [0:29] sb_1__1__0_chanx_right_out;
wire [0:29] sb_1__1__0_chany_bottom_out;
wire [0:29] sb_1__1__0_chany_top_out;
wire [0:29] sb_1__1__10_chanx_left_out;
wire [0:29] sb_1__1__10_chanx_right_out;
wire [0:29] sb_1__1__10_chany_bottom_out;
wire [0:29] sb_1__1__10_chany_top_out;
wire [0:29] sb_1__1__11_chanx_left_out;
wire [0:29] sb_1__1__11_chanx_right_out;
wire [0:29] sb_1__1__11_chany_bottom_out;
wire [0:29] sb_1__1__11_chany_top_out;
wire [0:29] sb_1__1__12_chanx_left_out;
wire [0:29] sb_1__1__12_chanx_right_out;
wire [0:29] sb_1__1__12_chany_bottom_out;
wire [0:29] sb_1__1__12_chany_top_out;
wire [0:29] sb_1__1__13_chanx_left_out;
wire [0:29] sb_1__1__13_chanx_right_out;
wire [0:29] sb_1__1__13_chany_bottom_out;
wire [0:29] sb_1__1__13_chany_top_out;
wire [0:29] sb_1__1__14_chanx_left_out;
wire [0:29] sb_1__1__14_chanx_right_out;
wire [0:29] sb_1__1__14_chany_bottom_out;
wire [0:29] sb_1__1__14_chany_top_out;
wire [0:29] sb_1__1__15_chanx_left_out;
wire [0:29] sb_1__1__15_chanx_right_out;
wire [0:29] sb_1__1__15_chany_bottom_out;
wire [0:29] sb_1__1__15_chany_top_out;
wire [0:29] sb_1__1__16_chanx_left_out;
wire [0:29] sb_1__1__16_chanx_right_out;
wire [0:29] sb_1__1__16_chany_bottom_out;
wire [0:29] sb_1__1__16_chany_top_out;
wire [0:29] sb_1__1__17_chanx_left_out;
wire [0:29] sb_1__1__17_chanx_right_out;
wire [0:29] sb_1__1__17_chany_bottom_out;
wire [0:29] sb_1__1__17_chany_top_out;
wire [0:29] sb_1__1__18_chanx_left_out;
wire [0:29] sb_1__1__18_chanx_right_out;
wire [0:29] sb_1__1__18_chany_bottom_out;
wire [0:29] sb_1__1__18_chany_top_out;
wire [0:29] sb_1__1__19_chanx_left_out;
wire [0:29] sb_1__1__19_chanx_right_out;
wire [0:29] sb_1__1__19_chany_bottom_out;
wire [0:29] sb_1__1__19_chany_top_out;
wire [0:29] sb_1__1__1_chanx_left_out;
wire [0:29] sb_1__1__1_chanx_right_out;
wire [0:29] sb_1__1__1_chany_bottom_out;
wire [0:29] sb_1__1__1_chany_top_out;
wire [0:29] sb_1__1__20_chanx_left_out;
wire [0:29] sb_1__1__20_chanx_right_out;
wire [0:29] sb_1__1__20_chany_bottom_out;
wire [0:29] sb_1__1__20_chany_top_out;
wire [0:29] sb_1__1__21_chanx_left_out;
wire [0:29] sb_1__1__21_chanx_right_out;
wire [0:29] sb_1__1__21_chany_bottom_out;
wire [0:29] sb_1__1__21_chany_top_out;
wire [0:29] sb_1__1__22_chanx_left_out;
wire [0:29] sb_1__1__22_chanx_right_out;
wire [0:29] sb_1__1__22_chany_bottom_out;
wire [0:29] sb_1__1__22_chany_top_out;
wire [0:29] sb_1__1__23_chanx_left_out;
wire [0:29] sb_1__1__23_chanx_right_out;
wire [0:29] sb_1__1__23_chany_bottom_out;
wire [0:29] sb_1__1__23_chany_top_out;
wire [0:29] sb_1__1__24_chanx_left_out;
wire [0:29] sb_1__1__24_chanx_right_out;
wire [0:29] sb_1__1__24_chany_bottom_out;
wire [0:29] sb_1__1__24_chany_top_out;
wire [0:29] sb_1__1__25_chanx_left_out;
wire [0:29] sb_1__1__25_chanx_right_out;
wire [0:29] sb_1__1__25_chany_bottom_out;
wire [0:29] sb_1__1__25_chany_top_out;
wire [0:29] sb_1__1__26_chanx_left_out;
wire [0:29] sb_1__1__26_chanx_right_out;
wire [0:29] sb_1__1__26_chany_bottom_out;
wire [0:29] sb_1__1__26_chany_top_out;
wire [0:29] sb_1__1__27_chanx_left_out;
wire [0:29] sb_1__1__27_chanx_right_out;
wire [0:29] sb_1__1__27_chany_bottom_out;
wire [0:29] sb_1__1__27_chany_top_out;
wire [0:29] sb_1__1__28_chanx_left_out;
wire [0:29] sb_1__1__28_chanx_right_out;
wire [0:29] sb_1__1__28_chany_bottom_out;
wire [0:29] sb_1__1__28_chany_top_out;
wire [0:29] sb_1__1__29_chanx_left_out;
wire [0:29] sb_1__1__29_chanx_right_out;
wire [0:29] sb_1__1__29_chany_bottom_out;
wire [0:29] sb_1__1__29_chany_top_out;
wire [0:29] sb_1__1__2_chanx_left_out;
wire [0:29] sb_1__1__2_chanx_right_out;
wire [0:29] sb_1__1__2_chany_bottom_out;
wire [0:29] sb_1__1__2_chany_top_out;
wire [0:29] sb_1__1__30_chanx_left_out;
wire [0:29] sb_1__1__30_chanx_right_out;
wire [0:29] sb_1__1__30_chany_bottom_out;
wire [0:29] sb_1__1__30_chany_top_out;
wire [0:29] sb_1__1__31_chanx_left_out;
wire [0:29] sb_1__1__31_chanx_right_out;
wire [0:29] sb_1__1__31_chany_bottom_out;
wire [0:29] sb_1__1__31_chany_top_out;
wire [0:29] sb_1__1__32_chanx_left_out;
wire [0:29] sb_1__1__32_chanx_right_out;
wire [0:29] sb_1__1__32_chany_bottom_out;
wire [0:29] sb_1__1__32_chany_top_out;
wire [0:29] sb_1__1__33_chanx_left_out;
wire [0:29] sb_1__1__33_chanx_right_out;
wire [0:29] sb_1__1__33_chany_bottom_out;
wire [0:29] sb_1__1__33_chany_top_out;
wire [0:29] sb_1__1__34_chanx_left_out;
wire [0:29] sb_1__1__34_chanx_right_out;
wire [0:29] sb_1__1__34_chany_bottom_out;
wire [0:29] sb_1__1__34_chany_top_out;
wire [0:29] sb_1__1__35_chanx_left_out;
wire [0:29] sb_1__1__35_chanx_right_out;
wire [0:29] sb_1__1__35_chany_bottom_out;
wire [0:29] sb_1__1__35_chany_top_out;
wire [0:29] sb_1__1__36_chanx_left_out;
wire [0:29] sb_1__1__36_chanx_right_out;
wire [0:29] sb_1__1__36_chany_bottom_out;
wire [0:29] sb_1__1__36_chany_top_out;
wire [0:29] sb_1__1__37_chanx_left_out;
wire [0:29] sb_1__1__37_chanx_right_out;
wire [0:29] sb_1__1__37_chany_bottom_out;
wire [0:29] sb_1__1__37_chany_top_out;
wire [0:29] sb_1__1__38_chanx_left_out;
wire [0:29] sb_1__1__38_chanx_right_out;
wire [0:29] sb_1__1__38_chany_bottom_out;
wire [0:29] sb_1__1__38_chany_top_out;
wire [0:29] sb_1__1__39_chanx_left_out;
wire [0:29] sb_1__1__39_chanx_right_out;
wire [0:29] sb_1__1__39_chany_bottom_out;
wire [0:29] sb_1__1__39_chany_top_out;
wire [0:29] sb_1__1__3_chanx_left_out;
wire [0:29] sb_1__1__3_chanx_right_out;
wire [0:29] sb_1__1__3_chany_bottom_out;
wire [0:29] sb_1__1__3_chany_top_out;
wire [0:29] sb_1__1__40_chanx_left_out;
wire [0:29] sb_1__1__40_chanx_right_out;
wire [0:29] sb_1__1__40_chany_bottom_out;
wire [0:29] sb_1__1__40_chany_top_out;
wire [0:29] sb_1__1__41_chanx_left_out;
wire [0:29] sb_1__1__41_chanx_right_out;
wire [0:29] sb_1__1__41_chany_bottom_out;
wire [0:29] sb_1__1__41_chany_top_out;
wire [0:29] sb_1__1__42_chanx_left_out;
wire [0:29] sb_1__1__42_chanx_right_out;
wire [0:29] sb_1__1__42_chany_bottom_out;
wire [0:29] sb_1__1__42_chany_top_out;
wire [0:29] sb_1__1__43_chanx_left_out;
wire [0:29] sb_1__1__43_chanx_right_out;
wire [0:29] sb_1__1__43_chany_bottom_out;
wire [0:29] sb_1__1__43_chany_top_out;
wire [0:29] sb_1__1__44_chanx_left_out;
wire [0:29] sb_1__1__44_chanx_right_out;
wire [0:29] sb_1__1__44_chany_bottom_out;
wire [0:29] sb_1__1__44_chany_top_out;
wire [0:29] sb_1__1__45_chanx_left_out;
wire [0:29] sb_1__1__45_chanx_right_out;
wire [0:29] sb_1__1__45_chany_bottom_out;
wire [0:29] sb_1__1__45_chany_top_out;
wire [0:29] sb_1__1__46_chanx_left_out;
wire [0:29] sb_1__1__46_chanx_right_out;
wire [0:29] sb_1__1__46_chany_bottom_out;
wire [0:29] sb_1__1__46_chany_top_out;
wire [0:29] sb_1__1__47_chanx_left_out;
wire [0:29] sb_1__1__47_chanx_right_out;
wire [0:29] sb_1__1__47_chany_bottom_out;
wire [0:29] sb_1__1__47_chany_top_out;
wire [0:29] sb_1__1__48_chanx_left_out;
wire [0:29] sb_1__1__48_chanx_right_out;
wire [0:29] sb_1__1__48_chany_bottom_out;
wire [0:29] sb_1__1__48_chany_top_out;
wire [0:29] sb_1__1__4_chanx_left_out;
wire [0:29] sb_1__1__4_chanx_right_out;
wire [0:29] sb_1__1__4_chany_bottom_out;
wire [0:29] sb_1__1__4_chany_top_out;
wire [0:29] sb_1__1__5_chanx_left_out;
wire [0:29] sb_1__1__5_chanx_right_out;
wire [0:29] sb_1__1__5_chany_bottom_out;
wire [0:29] sb_1__1__5_chany_top_out;
wire [0:29] sb_1__1__6_chanx_left_out;
wire [0:29] sb_1__1__6_chanx_right_out;
wire [0:29] sb_1__1__6_chany_bottom_out;
wire [0:29] sb_1__1__6_chany_top_out;
wire [0:29] sb_1__1__7_chanx_left_out;
wire [0:29] sb_1__1__7_chanx_right_out;
wire [0:29] sb_1__1__7_chany_bottom_out;
wire [0:29] sb_1__1__7_chany_top_out;
wire [0:29] sb_1__1__8_chanx_left_out;
wire [0:29] sb_1__1__8_chanx_right_out;
wire [0:29] sb_1__1__8_chany_bottom_out;
wire [0:29] sb_1__1__8_chany_top_out;
wire [0:29] sb_1__1__9_chanx_left_out;
wire [0:29] sb_1__1__9_chanx_right_out;
wire [0:29] sb_1__1__9_chany_bottom_out;
wire [0:29] sb_1__1__9_chany_top_out;
wire [0:29] sb_1__8__0_chanx_left_out;
wire [0:29] sb_1__8__0_chanx_right_out;
wire [0:29] sb_1__8__0_chany_bottom_out;
wire [0:29] sb_1__8__1_chanx_left_out;
wire [0:29] sb_1__8__1_chanx_right_out;
wire [0:29] sb_1__8__1_chany_bottom_out;
wire [0:29] sb_1__8__2_chanx_left_out;
wire [0:29] sb_1__8__2_chanx_right_out;
wire [0:29] sb_1__8__2_chany_bottom_out;
wire [0:29] sb_1__8__3_chanx_left_out;
wire [0:29] sb_1__8__3_chanx_right_out;
wire [0:29] sb_1__8__3_chany_bottom_out;
wire [0:29] sb_1__8__4_chanx_left_out;
wire [0:29] sb_1__8__4_chanx_right_out;
wire [0:29] sb_1__8__4_chany_bottom_out;
wire [0:29] sb_1__8__5_chanx_left_out;
wire [0:29] sb_1__8__5_chanx_right_out;
wire [0:29] sb_1__8__5_chany_bottom_out;
wire [0:29] sb_1__8__6_chanx_left_out;
wire [0:29] sb_1__8__6_chanx_right_out;
wire [0:29] sb_1__8__6_chany_bottom_out;
wire [0:29] sb_8__0__0_chanx_left_out;
wire [0:29] sb_8__0__0_chany_top_out;
wire [0:29] sb_8__1__0_chanx_left_out;
wire [0:29] sb_8__1__0_chany_bottom_out;
wire [0:29] sb_8__1__0_chany_top_out;
wire [0:29] sb_8__1__1_chanx_left_out;
wire [0:29] sb_8__1__1_chany_bottom_out;
wire [0:29] sb_8__1__1_chany_top_out;
wire [0:29] sb_8__1__2_chanx_left_out;
wire [0:29] sb_8__1__2_chany_bottom_out;
wire [0:29] sb_8__1__2_chany_top_out;
wire [0:29] sb_8__1__3_chanx_left_out;
wire [0:29] sb_8__1__3_chany_bottom_out;
wire [0:29] sb_8__1__3_chany_top_out;
wire [0:29] sb_8__1__4_chanx_left_out;
wire [0:29] sb_8__1__4_chany_bottom_out;
wire [0:29] sb_8__1__4_chany_top_out;
wire [0:29] sb_8__1__5_chanx_left_out;
wire [0:29] sb_8__1__5_chany_bottom_out;
wire [0:29] sb_8__1__5_chany_top_out;
wire [0:29] sb_8__1__6_chanx_left_out;
wire [0:29] sb_8__1__6_chany_bottom_out;
wire [0:29] sb_8__1__6_chany_top_out;
wire [0:29] sb_8__8__0_chanx_left_out;
wire [0:29] sb_8__8__0_chany_bottom_out;

// ----- BEGIN Local short connections -----
// ----- END Local short connections -----
// ----- BEGIN Local output short connections -----
// ----- END Local output short connections -----

	grid_io_top_top grid_io_top_top_1__9_ (
		.isol_n(isol_n),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[0:3]),
		.gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[0:3]),
		.gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[0:3]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__8__0_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__8__0_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__8__0_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__8__0_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.ccff_head(cbx_1__8__0_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_top_0_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_top_0_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_top_0_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.ccff_tail(grid_io_top_top_0_ccff_tail));

	grid_io_top_top grid_io_top_top_2__9_ (
		.isol_n(isol_n),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[4:7]),
		.gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[4:7]),
		.gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[4:7]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__8__1_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__8__1_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__8__1_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__8__1_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.ccff_head(cbx_1__8__1_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_top_1_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_top_1_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_top_1_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.ccff_tail(grid_io_top_top_1_ccff_tail));

	grid_io_top_top grid_io_top_top_3__9_ (
		.isol_n(isol_n),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[8:11]),
		.gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[8:11]),
		.gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[8:11]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__8__2_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__8__2_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__8__2_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__8__2_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.ccff_head(cbx_1__8__2_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_top_2_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_top_2_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_top_2_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.ccff_tail(grid_io_top_top_2_ccff_tail));

	grid_io_top_top grid_io_top_top_4__9_ (
		.isol_n(isol_n),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[12:15]),
		.gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[12:15]),
		.gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[12:15]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__8__3_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__8__3_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__8__3_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__8__3_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.ccff_head(cbx_1__8__3_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_top_3_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_top_3_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_top_3_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.ccff_tail(grid_io_top_top_3_ccff_tail));

	grid_io_top_top grid_io_top_top_5__9_ (
		.isol_n(isol_n),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[16:19]),
		.gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[16:19]),
		.gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[16:19]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__8__4_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__8__4_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__8__4_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__8__4_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.ccff_head(cbx_1__8__4_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_4_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_top_4_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_top_4_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_top_4_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.ccff_tail(grid_io_top_top_4_ccff_tail));

	grid_io_top_top grid_io_top_top_6__9_ (
		.isol_n(isol_n),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[20:23]),
		.gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[20:23]),
		.gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[20:23]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__8__5_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__8__5_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__8__5_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__8__5_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.ccff_head(cbx_1__8__5_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_5_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_top_5_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_top_5_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_top_5_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.ccff_tail(grid_io_top_top_5_ccff_tail));

	grid_io_top_top grid_io_top_top_7__9_ (
		.isol_n(isol_n),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[24:27]),
		.gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[24:27]),
		.gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[24:27]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__8__6_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__8__6_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__8__6_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__8__6_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.ccff_head(cbx_1__8__6_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_6_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_top_6_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_top_6_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_top_6_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.ccff_tail(grid_io_top_top_6_ccff_tail));

	grid_io_top_top grid_io_top_top_8__9_ (
		.isol_n(isol_n),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[28:31]),
		.gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[28:31]),
		.gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[28:31]),
		.bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__8__7_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__8__7_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__8__7_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__8__7_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.ccff_head(cbx_1__8__7_ccff_tail),
		.bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_7_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_top_7_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_top_7_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_top_7_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.ccff_tail(grid_io_top_top_7_ccff_tail));

	grid_io_right_right grid_io_right_right_9__8_ (
		.isol_n(isol_n),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[32:35]),
		.gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[32:35]),
		.gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[32:35]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_8__1__7_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_8__1__7_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_8__1__7_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_8__1__7_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.ccff_head(grid_io_right_right_1_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_right_0_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_right_0_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_right_0_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.ccff_tail(grid_io_right_right_0_ccff_tail));

	grid_io_right_right grid_io_right_right_9__7_ (
		.isol_n(isol_n),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[36:39]),
		.gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[36:39]),
		.gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[36:39]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_8__1__6_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_8__1__6_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_8__1__6_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_8__1__6_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.ccff_head(grid_io_right_right_2_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_right_1_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_right_1_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_right_1_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.ccff_tail(grid_io_right_right_1_ccff_tail));

	grid_io_right_right grid_io_right_right_9__6_ (
		.isol_n(isol_n),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[40:43]),
		.gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[40:43]),
		.gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[40:43]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_8__1__5_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_8__1__5_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_8__1__5_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_8__1__5_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.ccff_head(grid_io_right_right_3_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_right_2_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_right_2_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_right_2_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.ccff_tail(grid_io_right_right_2_ccff_tail));

	grid_io_right_right grid_io_right_right_9__5_ (
		.isol_n(isol_n),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[44:47]),
		.gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[44:47]),
		.gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[44:47]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_8__1__4_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_8__1__4_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_8__1__4_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_8__1__4_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.ccff_head(grid_io_right_right_4_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_3_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_right_3_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_right_3_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_right_3_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.ccff_tail(grid_io_right_right_3_ccff_tail));

	grid_io_right_right grid_io_right_right_9__4_ (
		.isol_n(isol_n),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[48:51]),
		.gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[48:51]),
		.gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[48:51]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_8__1__3_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_8__1__3_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_8__1__3_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_8__1__3_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.ccff_head(grid_io_right_right_5_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_4_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_right_4_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_right_4_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_right_4_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.ccff_tail(grid_io_right_right_4_ccff_tail));

	grid_io_right_right grid_io_right_right_9__3_ (
		.isol_n(isol_n),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[52:55]),
		.gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[52:55]),
		.gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[52:55]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_8__1__2_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_8__1__2_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_8__1__2_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_8__1__2_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.ccff_head(grid_io_right_right_6_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_5_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_right_5_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_right_5_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_right_5_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.ccff_tail(grid_io_right_right_5_ccff_tail));

	grid_io_right_right grid_io_right_right_9__2_ (
		.isol_n(isol_n),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[56:59]),
		.gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[56:59]),
		.gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[56:59]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_8__1__1_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_8__1__1_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_8__1__1_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_8__1__1_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.ccff_head(grid_io_right_right_7_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_6_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_right_6_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_right_6_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_right_6_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.ccff_tail(grid_io_right_right_6_ccff_tail));

	grid_io_right_right grid_io_right_right_9__1_ (
		.isol_n(isol_n),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[60:63]),
		.gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[60:63]),
		.gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[60:63]),
		.left_width_0_height_0_subtile_0__pin_outpad_0_(cby_8__1__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_width_0_height_0_subtile_1__pin_outpad_0_(cby_8__1__0_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_width_0_height_0_subtile_2__pin_outpad_0_(cby_8__1__0_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_width_0_height_0_subtile_3__pin_outpad_0_(cby_8__1__0_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.ccff_head(grid_io_bottom_bottom_0_ccff_tail),
		.left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_7_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_right_7_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_right_7_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_right_7_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.ccff_tail(grid_io_right_right_7_ccff_tail));

	grid_io_bottom_bottom grid_io_bottom_bottom_8__0_ (
		.isol_n(isol_n),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[64:67]),
		.gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[64:67]),
		.gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[64:67]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.ccff_head(grid_io_bottom_bottom_1_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_bottom_0_ccff_tail));

	grid_io_bottom_bottom grid_io_bottom_bottom_7__0_ (
		.isol_n(isol_n),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[68:71]),
		.gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[68:71]),
		.gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[68:71]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.ccff_head(grid_io_bottom_bottom_2_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_bottom_1_ccff_tail));

	grid_io_bottom_bottom grid_io_bottom_bottom_6__0_ (
		.isol_n(isol_n),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[72:75]),
		.gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[72:75]),
		.gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[72:75]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.ccff_head(grid_io_bottom_bottom_3_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_bottom_2_ccff_tail));

	grid_io_bottom_bottom grid_io_bottom_bottom_5__0_ (
		.isol_n(isol_n),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[76:79]),
		.gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[76:79]),
		.gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[76:79]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.ccff_head(grid_io_bottom_bottom_4_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_bottom_3_ccff_tail));

	grid_io_bottom_bottom grid_io_bottom_bottom_4__0_ (
		.isol_n(isol_n),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[80:83]),
		.gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[80:83]),
		.gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[80:83]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.ccff_head(grid_io_bottom_bottom_5_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_bottom_4_ccff_tail));

	grid_io_bottom_bottom grid_io_bottom_bottom_3__0_ (
		.isol_n(isol_n),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[84:87]),
		.gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[84:87]),
		.gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[84:87]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.ccff_head(grid_io_bottom_bottom_6_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_bottom_5_ccff_tail));

	grid_io_bottom_bottom grid_io_bottom_bottom_2__0_ (
		.isol_n(isol_n),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[88:91]),
		.gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[88:91]),
		.gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[88:91]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.ccff_head(grid_io_bottom_bottom_7_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_bottom_6_ccff_tail));

	grid_io_bottom_bottom grid_io_bottom_bottom_1__0_ (
		.isol_n(isol_n),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[92:95]),
		.gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[92:95]),
		.gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[92:95]),
		.top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.ccff_head(ccff_head),
		.top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.ccff_tail(grid_io_bottom_bottom_7_ccff_tail));

	grid_io_left_left grid_io_left_left_0__1_ (
		.isol_n(isol_n),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[96:99]),
		.gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[96:99]),
		.gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[96:99]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.ccff_head(cby_0__1__0_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_left_0_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_left_0_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_left_0_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.ccff_tail(grid_io_left_left_0_ccff_tail));

	grid_io_left_left grid_io_left_left_0__2_ (
		.isol_n(isol_n),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[100:103]),
		.gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[100:103]),
		.gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[100:103]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.ccff_head(cby_0__1__1_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_left_1_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_left_1_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_left_1_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.ccff_tail(grid_io_left_left_1_ccff_tail));

	grid_io_left_left grid_io_left_left_0__3_ (
		.isol_n(isol_n),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[104:107]),
		.gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[104:107]),
		.gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[104:107]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.ccff_head(cby_0__1__2_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_left_2_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_left_2_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_left_2_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.ccff_tail(grid_io_left_left_2_ccff_tail));

	grid_io_left_left grid_io_left_left_0__4_ (
		.isol_n(isol_n),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[108:111]),
		.gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[108:111]),
		.gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[108:111]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.ccff_head(cby_0__1__3_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_3_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_left_3_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_left_3_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_left_3_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.ccff_tail(grid_io_left_left_3_ccff_tail));

	grid_io_left_left grid_io_left_left_0__5_ (
		.isol_n(isol_n),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[112:115]),
		.gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[112:115]),
		.gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[112:115]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.ccff_head(cby_0__1__4_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_4_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_left_4_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_left_4_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_left_4_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.ccff_tail(grid_io_left_left_4_ccff_tail));

	grid_io_left_left grid_io_left_left_0__6_ (
		.isol_n(isol_n),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[116:119]),
		.gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[116:119]),
		.gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[116:119]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__5_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__5_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__5_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__5_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.ccff_head(cby_0__1__5_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_5_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_left_5_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_left_5_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_left_5_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.ccff_tail(grid_io_left_left_5_ccff_tail));

	grid_io_left_left grid_io_left_left_0__7_ (
		.isol_n(isol_n),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[120:123]),
		.gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[120:123]),
		.gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[120:123]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__6_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__6_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__6_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__6_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.ccff_head(cby_0__1__6_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_6_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_left_6_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_left_6_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_left_6_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.ccff_tail(grid_io_left_left_6_ccff_tail));

	grid_io_left_left grid_io_left_left_0__8_ (
		.isol_n(isol_n),
		.pReset(pReset),
		.prog_clk(prog_clk),
		.gfpga_pad_io_soc_in(gfpga_pad_io_soc_in[124:127]),
		.gfpga_pad_io_soc_out(gfpga_pad_io_soc_out[124:127]),
		.gfpga_pad_io_soc_dir(gfpga_pad_io_soc_dir[124:127]),
		.right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__7_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__7_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__7_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__7_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.ccff_head(cby_0__1__7_ccff_tail),
		.right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_7_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_left_7_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_left_7_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_left_7_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.ccff_tail(grid_io_left_left_7_ccff_tail));

	grid_clb grid_clb_1__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_56_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_112_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_0_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__0_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_1__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_0_ccff_tail));

	grid_clb grid_clb_1__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_57_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_113_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_1_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__1_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_1_ccff_tail));

	grid_clb grid_clb_1__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_58_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_114_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_2_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__2_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_2_ccff_tail));

	grid_clb grid_clb_1__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_59_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_115_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_3_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__3_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_3_ccff_tail));

	grid_clb grid_clb_1__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_60_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_116_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_4_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__4_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_4_ccff_tail));

	grid_clb grid_clb_1__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_61_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_117_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_5_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__5_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_5_ccff_tail));

	grid_clb grid_clb_1__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_62_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_118_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_6_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__6_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_6_ccff_tail));

	grid_clb grid_clb_1__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__8__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__8__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__8__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__8__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__8__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__8__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__8__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__8__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__8__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__8__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__8__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__8__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__8__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__8__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__8__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__8__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_1__8__undriven_top_width_0_height_0_subtile_0__pin_reg_in_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(grid_clb_1__8__undriven_top_width_0_height_0_subtile_0__pin_sc_in_0_),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_1__8__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__7_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(ccff_tail));

	grid_clb grid_clb_2__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_63_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_119_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_7_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__8_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_8_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_2__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_8_ccff_tail));

	grid_clb grid_clb_2__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_64_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_120_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_8_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__9_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_9_ccff_tail));

	grid_clb grid_clb_2__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_65_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_121_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_9_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__10_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_10_ccff_tail));

	grid_clb grid_clb_2__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_66_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_122_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_10_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__11_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_11_ccff_tail));

	grid_clb grid_clb_2__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_67_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_123_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_11_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__12_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_12_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_12_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_12_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_12_ccff_tail));

	grid_clb grid_clb_2__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_68_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_124_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_12_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__13_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_13_ccff_tail));

	grid_clb grid_clb_2__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_69_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_125_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_13_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__14_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_14_ccff_tail));

	grid_clb grid_clb_2__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__8__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__8__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__8__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__8__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__8__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__8__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__8__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__8__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__8__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__8__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__8__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__8__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__8__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__8__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__8__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__8__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_2__8__undriven_top_width_0_height_0_subtile_0__pin_reg_in_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_168_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_2__8__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__15_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_15_ccff_tail));

	grid_clb grid_clb_3__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_70_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_126_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_14_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__16_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_16_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_3__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_16_ccff_tail));

	grid_clb grid_clb_3__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_71_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_127_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_15_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__17_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_17_ccff_tail));

	grid_clb grid_clb_3__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_72_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_128_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_16_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__18_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_18_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_18_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_18_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_18_ccff_tail));

	grid_clb grid_clb_3__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_73_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_129_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_17_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__19_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_19_ccff_tail));

	grid_clb grid_clb_3__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_74_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_130_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_18_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__20_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_20_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_20_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_20_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_20_ccff_tail));

	grid_clb grid_clb_3__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_75_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_131_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_19_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__21_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_21_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_21_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_21_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_21_ccff_tail));

	grid_clb grid_clb_3__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_76_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_132_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_20_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__22_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_22_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_22_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_22_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_22_ccff_tail));

	grid_clb grid_clb_3__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__8__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__8__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__8__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__8__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__8__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__8__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__8__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__8__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__8__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__8__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__8__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__8__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__8__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__8__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__8__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__8__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_3__8__undriven_top_width_0_height_0_subtile_0__pin_reg_in_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_169_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_3__8__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__23_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_23_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_23_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_23_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_23_ccff_tail));

	grid_clb grid_clb_4__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_77_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_133_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_21_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__24_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_24_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_4__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_24_ccff_tail));

	grid_clb grid_clb_4__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_78_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_134_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_22_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__25_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_25_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_25_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_25_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_25_ccff_tail));

	grid_clb grid_clb_4__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_79_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_135_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_23_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__26_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_26_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_26_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_26_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_26_ccff_tail));

	grid_clb grid_clb_4__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_80_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_136_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_24_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__27_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_27_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_27_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_27_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_27_ccff_tail));

	grid_clb grid_clb_4__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_81_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_137_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_25_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__28_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_28_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_28_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_28_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_28_ccff_tail));

	grid_clb grid_clb_4__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_82_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_138_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_26_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__29_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_29_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_29_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_29_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_29_ccff_tail));

	grid_clb grid_clb_4__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_83_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_139_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_27_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__30_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_30_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_30_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_30_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_30_ccff_tail));

	grid_clb grid_clb_4__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__8__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__8__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__8__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__8__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__8__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__8__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__8__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__8__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__8__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__8__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__8__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__8__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__8__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__8__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__8__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__8__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_4__8__undriven_top_width_0_height_0_subtile_0__pin_reg_in_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_170_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_4__8__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__31_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_31_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_31_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_31_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_31_ccff_tail));

	grid_clb grid_clb_5__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_84_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_140_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_28_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__32_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_32_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_5__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_32_ccff_tail));

	grid_clb grid_clb_5__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_85_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_141_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_29_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__33_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_33_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_33_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_33_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_33_ccff_tail));

	grid_clb grid_clb_5__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_86_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_142_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_30_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__34_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_34_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_34_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_34_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_34_ccff_tail));

	grid_clb grid_clb_5__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_87_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_143_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_31_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__35_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_35_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_35_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_35_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_35_ccff_tail));

	grid_clb grid_clb_5__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_88_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_144_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_32_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__36_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_36_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_36_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_36_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_36_ccff_tail));

	grid_clb grid_clb_5__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_89_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_145_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_33_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__37_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_37_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_37_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_37_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_37_ccff_tail));

	grid_clb grid_clb_5__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_90_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_146_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_34_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__38_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_38_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_38_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_38_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_38_ccff_tail));

	grid_clb grid_clb_5__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__8__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__8__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__8__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__8__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__8__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__8__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__8__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__8__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__8__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__8__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__8__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__8__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__8__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__8__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__8__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__8__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_5__8__undriven_top_width_0_height_0_subtile_0__pin_reg_in_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_171_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_5__8__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__39_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_39_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_39_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_39_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_39_ccff_tail));

	grid_clb grid_clb_6__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_91_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_147_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_35_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__40_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_6__1__undriven_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_40_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_6__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_40_ccff_tail));

	grid_clb grid_clb_6__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_92_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_148_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_36_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__41_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_41_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_41_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_41_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_41_ccff_tail));

	grid_clb grid_clb_6__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_93_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_149_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_37_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__42_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_42_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_42_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_42_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_42_ccff_tail));

	grid_clb grid_clb_6__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_94_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_150_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_38_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__43_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_43_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_43_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_43_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_43_ccff_tail));

	grid_clb grid_clb_6__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_95_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_151_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_39_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__44_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_44_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_44_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_44_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_44_ccff_tail));

	grid_clb grid_clb_6__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_96_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_152_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_40_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__45_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_45_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_45_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_45_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_45_ccff_tail));

	grid_clb grid_clb_6__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_97_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_153_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_41_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__46_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_46_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_46_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_46_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_46_ccff_tail));

	grid_clb grid_clb_6__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__8__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__8__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__8__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__8__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__8__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__8__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__8__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__8__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__8__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__8__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__8__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__8__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__8__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__8__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__8__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__8__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_6__8__undriven_top_width_0_height_0_subtile_0__pin_reg_in_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_172_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_6__8__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__47_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_47_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_47_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_47_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_47_ccff_tail));

	grid_clb grid_clb_7__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_98_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_154_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_42_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__48_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_48_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_7__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_48_ccff_tail));

	grid_clb grid_clb_7__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_99_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_155_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_43_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__49_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_49_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_49_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_49_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_49_ccff_tail));

	grid_clb grid_clb_7__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_100_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_156_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_44_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__50_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_50_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_50_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_50_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_50_ccff_tail));

	grid_clb grid_clb_7__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_101_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_157_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_45_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__51_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_51_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_51_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_51_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_51_ccff_tail));

	grid_clb grid_clb_7__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_102_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_158_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_46_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__52_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_52_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_52_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_52_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_52_ccff_tail));

	grid_clb grid_clb_7__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_103_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_159_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_47_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__53_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_53_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_53_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_53_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_53_ccff_tail));

	grid_clb grid_clb_7__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_104_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_160_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_48_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__54_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_54_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_54_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_54_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_54_ccff_tail));

	grid_clb grid_clb_7__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__8__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__8__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__8__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__8__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__8__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__8__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__8__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__8__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__8__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__8__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__8__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__8__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__8__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__8__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__8__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__8__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_7__8__undriven_top_width_0_height_0_subtile_0__pin_reg_in_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_173_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_7__8__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_1__1__55_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_55_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_55_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_55_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_55_ccff_tail));

	grid_clb grid_clb_8__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_105_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_161_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_49_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_8__1__0_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_8__1__undriven_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_8__1__undriven_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_8__1__undriven_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_56_ccff_tail));

	grid_clb grid_clb_8__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_106_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_162_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_50_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_8__1__1_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_57_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_57_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_57_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_57_ccff_tail));

	grid_clb grid_clb_8__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_107_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_163_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_51_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_8__1__2_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_58_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_58_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_58_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_58_ccff_tail));

	grid_clb grid_clb_8__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_108_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_164_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_52_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_8__1__3_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_59_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_59_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_59_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_59_ccff_tail));

	grid_clb grid_clb_8__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_109_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_165_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_53_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_8__1__4_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_60_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_60_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_60_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_60_ccff_tail));

	grid_clb grid_clb_8__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_110_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_166_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_54_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_8__1__5_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_61_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_61_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_61_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_61_ccff_tail));

	grid_clb grid_clb_8__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(direct_interc_111_out),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_167_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(direct_interc_55_out),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_8__1__6_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_62_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_62_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_62_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_62_ccff_tail));

	grid_clb grid_clb_8__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.Test_en(Test_en),
		.top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__8__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__8__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__8__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__8__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__8__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__8__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__8__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__8__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__8__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__8__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__8__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__8__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__8__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__8__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__8__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__8__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.top_width_0_height_0_subtile_0__pin_reg_in_0_(grid_clb_8__8__undriven_top_width_0_height_0_subtile_0__pin_reg_in_0_),
		.top_width_0_height_0_subtile_0__pin_sc_in_0_(direct_interc_174_out),
		.top_width_0_height_0_subtile_0__pin_cin_0_(grid_clb_8__8__undriven_top_width_0_height_0_subtile_0__pin_cin_0_),
		.right_width_0_height_0_subtile_0__pin_I4_0_(cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.right_width_0_height_0_subtile_0__pin_I4_1_(cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.right_width_0_height_0_subtile_0__pin_I4i_0_(cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.right_width_0_height_0_subtile_0__pin_I4i_1_(cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.right_width_0_height_0_subtile_0__pin_I5_0_(cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.right_width_0_height_0_subtile_0__pin_I5_1_(cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.right_width_0_height_0_subtile_0__pin_I5i_0_(cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.right_width_0_height_0_subtile_0__pin_I5i_1_(cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.right_width_0_height_0_subtile_0__pin_I6_0_(cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.right_width_0_height_0_subtile_0__pin_I6_1_(cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.right_width_0_height_0_subtile_0__pin_I6i_0_(cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.right_width_0_height_0_subtile_0__pin_I6i_1_(cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.right_width_0_height_0_subtile_0__pin_I7_0_(cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.right_width_0_height_0_subtile_0__pin_I7_1_(cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.right_width_0_height_0_subtile_0__pin_I7i_0_(cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.right_width_0_height_0_subtile_0__pin_I7i_1_(cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.left_width_0_height_0_subtile_0__pin_reset_0_(reset),
		.left_width_0_height_0_subtile_0__pin_clk_0_(clk),
		.ccff_head(cby_8__1__7_ccff_tail),
		.top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_0_),
		.top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_1_),
		.top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_2_),
		.top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_3_),
		.top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_4_),
		.top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_5_),
		.top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_6_),
		.top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_7_),
		.right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_8_),
		.right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_9_),
		.right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_10_),
		.right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_11_),
		.right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_12_),
		.right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_13_),
		.right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_14_),
		.right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_15_),
		.bottom_width_0_height_0_subtile_0__pin_reg_out_0_(grid_clb_63_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_sc_out_0_(grid_clb_63_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.bottom_width_0_height_0_subtile_0__pin_cout_0_(grid_clb_63_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.ccff_tail(grid_clb_63_ccff_tail));

	sb_0__0_ sb_0__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__0_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_left_0_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_left_0_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_left_0_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.chanx_right_in(cbx_1__0__0_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.ccff_head(grid_io_left_left_1_ccff_tail),
		.chany_top_out(sb_0__0__0_chany_top_out[0:29]),
		.chanx_right_out(sb_0__0__0_chanx_right_out[0:29]),
		.ccff_tail(sb_0__0__0_ccff_tail));

	sb_0__1_ sb_0__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__1_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_left_1_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_left_1_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_left_1_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.chanx_right_in(cbx_1__1__0_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_0__1__0_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_0_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_left_0_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_left_0_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_left_0_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.ccff_head(grid_io_left_left_2_ccff_tail),
		.chany_top_out(sb_0__1__0_chany_top_out[0:29]),
		.chanx_right_out(sb_0__1__0_chanx_right_out[0:29]),
		.chany_bottom_out(sb_0__1__0_chany_bottom_out[0:29]),
		.ccff_tail(sb_0__1__0_ccff_tail));

	sb_0__1_ sb_0__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__2_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_left_2_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_left_2_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_left_2_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.chanx_right_in(cbx_1__1__1_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_0__1__1_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_1_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_left_1_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_left_1_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_left_1_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.ccff_head(grid_io_left_left_3_ccff_tail),
		.chany_top_out(sb_0__1__1_chany_top_out[0:29]),
		.chanx_right_out(sb_0__1__1_chanx_right_out[0:29]),
		.chany_bottom_out(sb_0__1__1_chany_bottom_out[0:29]),
		.ccff_tail(sb_0__1__1_ccff_tail));

	sb_0__1_ sb_0__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__3_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_3_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_left_3_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_left_3_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_left_3_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.chanx_right_in(cbx_1__1__2_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_0__1__2_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_2_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_left_2_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_left_2_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_left_2_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.ccff_head(grid_io_left_left_4_ccff_tail),
		.chany_top_out(sb_0__1__2_chany_top_out[0:29]),
		.chanx_right_out(sb_0__1__2_chanx_right_out[0:29]),
		.chany_bottom_out(sb_0__1__2_chany_bottom_out[0:29]),
		.ccff_tail(sb_0__1__2_ccff_tail));

	sb_0__1_ sb_0__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__4_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_4_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_left_4_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_left_4_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_left_4_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.chanx_right_in(cbx_1__1__3_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_0__1__3_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_3_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_left_3_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_left_3_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_left_3_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.ccff_head(grid_io_left_left_5_ccff_tail),
		.chany_top_out(sb_0__1__3_chany_top_out[0:29]),
		.chanx_right_out(sb_0__1__3_chanx_right_out[0:29]),
		.chany_bottom_out(sb_0__1__3_chany_bottom_out[0:29]),
		.ccff_tail(sb_0__1__3_ccff_tail));

	sb_0__1_ sb_0__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__5_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_5_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_left_5_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_left_5_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_left_5_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.chanx_right_in(cbx_1__1__4_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_0__1__4_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_4_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_left_4_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_left_4_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_left_4_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.ccff_head(grid_io_left_left_6_ccff_tail),
		.chany_top_out(sb_0__1__4_chany_top_out[0:29]),
		.chanx_right_out(sb_0__1__4_chanx_right_out[0:29]),
		.chany_bottom_out(sb_0__1__4_chany_bottom_out[0:29]),
		.ccff_tail(sb_0__1__4_ccff_tail));

	sb_0__1_ sb_0__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__6_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_6_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_left_6_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_left_6_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_left_6_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.chanx_right_in(cbx_1__1__5_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_0__1__5_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_5_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_left_5_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_left_5_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_left_5_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.ccff_head(grid_io_left_left_7_ccff_tail),
		.chany_top_out(sb_0__1__5_chany_top_out[0:29]),
		.chanx_right_out(sb_0__1__5_chanx_right_out[0:29]),
		.chany_bottom_out(sb_0__1__5_chany_bottom_out[0:29]),
		.ccff_tail(sb_0__1__5_ccff_tail));

	sb_0__1_ sb_0__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_0__1__7_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_7_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_left_7_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_left_7_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_left_7_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.chanx_right_in(cbx_1__1__6_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_0__1__6_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_6_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_left_6_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_left_6_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_left_6_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.ccff_head(sb_0__8__0_ccff_tail),
		.chany_top_out(sb_0__1__6_chany_top_out[0:29]),
		.chanx_right_out(sb_0__1__6_chanx_right_out[0:29]),
		.chany_bottom_out(sb_0__1__6_chany_bottom_out[0:29]),
		.ccff_tail(sb_0__1__6_ccff_tail));

	sb_0__8_ sb_0__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__8__0_chanx_left_out[0:29]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_top_0_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_top_0_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_top_0_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_0__1__7_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_left_left_7_right_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_left_left_7_right_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_left_left_7_right_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_left_left_7_right_width_0_height_0_subtile_3__pin_inpad_0_),
		.ccff_head(grid_io_top_top_0_ccff_tail),
		.chanx_right_out(sb_0__8__0_chanx_right_out[0:29]),
		.chany_bottom_out(sb_0__8__0_chany_bottom_out[0:29]),
		.ccff_tail(sb_0__8__0_ccff_tail));

	sb_1__0_ sb_1__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__0_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__0__1_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__0_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_7_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.ccff_head(grid_io_left_left_0_ccff_tail),
		.chany_top_out(sb_1__0__0_chany_top_out[0:29]),
		.chanx_right_out(sb_1__0__0_chanx_right_out[0:29]),
		.chanx_left_out(sb_1__0__0_chanx_left_out[0:29]),
		.ccff_tail(sb_1__0__0_ccff_tail));

	sb_1__0_ sb_2__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__8_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__0__2_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__1_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_6_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.ccff_head(grid_clb_0_ccff_tail),
		.chany_top_out(sb_1__0__1_chany_top_out[0:29]),
		.chanx_right_out(sb_1__0__1_chanx_right_out[0:29]),
		.chanx_left_out(sb_1__0__1_chanx_left_out[0:29]),
		.ccff_tail(sb_1__0__1_ccff_tail));

	sb_1__0_ sb_3__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__16_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__0__3_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__2_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_5_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.ccff_head(grid_clb_8_ccff_tail),
		.chany_top_out(sb_1__0__2_chany_top_out[0:29]),
		.chanx_right_out(sb_1__0__2_chanx_right_out[0:29]),
		.chanx_left_out(sb_1__0__2_chanx_left_out[0:29]),
		.ccff_tail(sb_1__0__2_ccff_tail));

	sb_1__0_ sb_4__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__24_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__0__4_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__3_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_4_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.ccff_head(grid_clb_16_ccff_tail),
		.chany_top_out(sb_1__0__3_chany_top_out[0:29]),
		.chanx_right_out(sb_1__0__3_chanx_right_out[0:29]),
		.chanx_left_out(sb_1__0__3_chanx_left_out[0:29]),
		.ccff_tail(sb_1__0__3_ccff_tail));

	sb_1__0_ sb_5__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__32_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__0__5_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__4_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_3_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.ccff_head(grid_clb_24_ccff_tail),
		.chany_top_out(sb_1__0__4_chany_top_out[0:29]),
		.chanx_right_out(sb_1__0__4_chanx_right_out[0:29]),
		.chanx_left_out(sb_1__0__4_chanx_left_out[0:29]),
		.ccff_tail(sb_1__0__4_ccff_tail));

	sb_1__0_ sb_6__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__40_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__0__6_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__5_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_2_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.ccff_head(grid_clb_32_ccff_tail),
		.chany_top_out(sb_1__0__5_chany_top_out[0:29]),
		.chanx_right_out(sb_1__0__5_chanx_right_out[0:29]),
		.chanx_left_out(sb_1__0__5_chanx_left_out[0:29]),
		.ccff_tail(sb_1__0__5_ccff_tail));

	sb_1__0_ sb_7__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__48_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__0__7_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__6_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_1_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.ccff_head(grid_clb_40_ccff_tail),
		.chany_top_out(sb_1__0__6_chany_top_out[0:29]),
		.chanx_right_out(sb_1__0__6_chanx_right_out[0:29]),
		.chanx_left_out(sb_1__0__6_chanx_left_out[0:29]),
		.ccff_tail(sb_1__0__6_ccff_tail));

	sb_1__1_ sb_1__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__1_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__7_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__0_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_0_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__0_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_0_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_9_ccff_tail),
		.chany_top_out(sb_1__1__0_chany_top_out[0:29]),
		.chanx_right_out(sb_1__1__0_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__1__0_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__1__0_chanx_left_out[0:29]),
		.ccff_tail(sb_1__1__0_ccff_tail));

	sb_1__1_ sb_1__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__2_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__8_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__1_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_1_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__1_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_1_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_1_ccff_tail),
		.chany_top_out(sb_1__1__1_chany_top_out[0:29]),
		.chanx_right_out(sb_1__1__1_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__1__1_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__1__1_chanx_left_out[0:29]),
		.ccff_tail(sb_1__1__1_ccff_tail));

	sb_1__1_ sb_1__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__3_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__9_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__2_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_2_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__2_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_2_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_11_ccff_tail),
		.chany_top_out(sb_1__1__2_chany_top_out[0:29]),
		.chanx_right_out(sb_1__1__2_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__1__2_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__1__2_chanx_left_out[0:29]),
		.ccff_tail(sb_1__1__2_ccff_tail));

	sb_1__1_ sb_1__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__4_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__10_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__3_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_3_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__3_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_3_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_3_ccff_tail),
		.chany_top_out(sb_1__1__3_chany_top_out[0:29]),
		.chanx_right_out(sb_1__1__3_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__1__3_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__1__3_chanx_left_out[0:29]),
		.ccff_tail(sb_1__1__3_ccff_tail));

	sb_1__1_ sb_1__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__5_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__11_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__4_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_4_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__4_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_4_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_13_ccff_tail),
		.chany_top_out(sb_1__1__4_chany_top_out[0:29]),
		.chanx_right_out(sb_1__1__4_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__1__4_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__1__4_chanx_left_out[0:29]),
		.ccff_tail(sb_1__1__4_ccff_tail));

	sb_1__1_ sb_1__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__6_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__12_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__5_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_5_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__5_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_5_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_5_ccff_tail),
		.chany_top_out(sb_1__1__5_chany_top_out[0:29]),
		.chanx_right_out(sb_1__1__5_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__1__5_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__1__5_chanx_left_out[0:29]),
		.ccff_tail(sb_1__1__5_ccff_tail));

	sb_1__1_ sb_1__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__7_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__13_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__6_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_6_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__6_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_6_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_15_ccff_tail),
		.chany_top_out(sb_1__1__6_chany_top_out[0:29]),
		.chanx_right_out(sb_1__1__6_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__1__6_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__1__6_chanx_left_out[0:29]),
		.ccff_tail(sb_1__1__6_ccff_tail));

	sb_1__1_ sb_2__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__9_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__14_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__8_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_8_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__7_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_8_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_17_ccff_tail),
		.chany_top_out(sb_1__1__7_chany_top_out[0:29]),
		.chanx_right_out(sb_1__1__7_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__1__7_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__1__7_chanx_left_out[0:29]),
		.ccff_tail(sb_1__1__7_ccff_tail));

	sb_1__1_ sb_2__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__10_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__15_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__9_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_9_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__8_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_9_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_2_ccff_tail),
		.chany_top_out(sb_1__1__8_chany_top_out[0:29]),
		.chanx_right_out(sb_1__1__8_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__1__8_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__1__8_chanx_left_out[0:29]),
		.ccff_tail(sb_1__1__8_ccff_tail));

	sb_1__1_ sb_2__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__11_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__16_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__10_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_10_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__9_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_10_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_19_ccff_tail),
		.chany_top_out(sb_1__1__9_chany_top_out[0:29]),
		.chanx_right_out(sb_1__1__9_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__1__9_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__1__9_chanx_left_out[0:29]),
		.ccff_tail(sb_1__1__9_ccff_tail));

	sb_1__1_ sb_2__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__12_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__17_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__11_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_11_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__10_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_11_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_4_ccff_tail),
		.chany_top_out(sb_1__1__10_chany_top_out[0:29]),
		.chanx_right_out(sb_1__1__10_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__1__10_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__1__10_chanx_left_out[0:29]),
		.ccff_tail(sb_1__1__10_ccff_tail));

	sb_1__1_ sb_2__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__13_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__18_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__12_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_12_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__11_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_12_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_21_ccff_tail),
		.chany_top_out(sb_1__1__11_chany_top_out[0:29]),
		.chanx_right_out(sb_1__1__11_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__1__11_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__1__11_chanx_left_out[0:29]),
		.ccff_tail(sb_1__1__11_ccff_tail));

	sb_1__1_ sb_2__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__14_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__19_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__13_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_13_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__12_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_13_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_6_ccff_tail),
		.chany_top_out(sb_1__1__12_chany_top_out[0:29]),
		.chanx_right_out(sb_1__1__12_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__1__12_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__1__12_chanx_left_out[0:29]),
		.ccff_tail(sb_1__1__12_ccff_tail));

	sb_1__1_ sb_2__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__15_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__20_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__14_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_14_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__13_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_14_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_23_ccff_tail),
		.chany_top_out(sb_1__1__13_chany_top_out[0:29]),
		.chanx_right_out(sb_1__1__13_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__1__13_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__1__13_chanx_left_out[0:29]),
		.ccff_tail(sb_1__1__13_ccff_tail));

	sb_1__1_ sb_3__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__17_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__21_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__16_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_16_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__14_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_16_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_25_ccff_tail),
		.chany_top_out(sb_1__1__14_chany_top_out[0:29]),
		.chanx_right_out(sb_1__1__14_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__1__14_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__1__14_chanx_left_out[0:29]),
		.ccff_tail(sb_1__1__14_ccff_tail));

	sb_1__1_ sb_3__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__18_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__22_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__17_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_17_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__15_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_17_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_10_ccff_tail),
		.chany_top_out(sb_1__1__15_chany_top_out[0:29]),
		.chanx_right_out(sb_1__1__15_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__1__15_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__1__15_chanx_left_out[0:29]),
		.ccff_tail(sb_1__1__15_ccff_tail));

	sb_1__1_ sb_3__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__19_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__23_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__18_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_18_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__16_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_18_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_27_ccff_tail),
		.chany_top_out(sb_1__1__16_chany_top_out[0:29]),
		.chanx_right_out(sb_1__1__16_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__1__16_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__1__16_chanx_left_out[0:29]),
		.ccff_tail(sb_1__1__16_ccff_tail));

	sb_1__1_ sb_3__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__20_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__24_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__19_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_19_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__17_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_19_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_12_ccff_tail),
		.chany_top_out(sb_1__1__17_chany_top_out[0:29]),
		.chanx_right_out(sb_1__1__17_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__1__17_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__1__17_chanx_left_out[0:29]),
		.ccff_tail(sb_1__1__17_ccff_tail));

	sb_1__1_ sb_3__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__21_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__25_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__20_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_20_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__18_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_20_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_29_ccff_tail),
		.chany_top_out(sb_1__1__18_chany_top_out[0:29]),
		.chanx_right_out(sb_1__1__18_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__1__18_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__1__18_chanx_left_out[0:29]),
		.ccff_tail(sb_1__1__18_ccff_tail));

	sb_1__1_ sb_3__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__22_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__26_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__21_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_21_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__19_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_21_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_14_ccff_tail),
		.chany_top_out(sb_1__1__19_chany_top_out[0:29]),
		.chanx_right_out(sb_1__1__19_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__1__19_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__1__19_chanx_left_out[0:29]),
		.ccff_tail(sb_1__1__19_ccff_tail));

	sb_1__1_ sb_3__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__23_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__27_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__22_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_22_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__20_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_22_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_31_ccff_tail),
		.chany_top_out(sb_1__1__20_chany_top_out[0:29]),
		.chanx_right_out(sb_1__1__20_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__1__20_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__1__20_chanx_left_out[0:29]),
		.ccff_tail(sb_1__1__20_ccff_tail));

	sb_1__1_ sb_4__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__25_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__28_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__24_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_24_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__21_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_24_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_33_ccff_tail),
		.chany_top_out(sb_1__1__21_chany_top_out[0:29]),
		.chanx_right_out(sb_1__1__21_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__1__21_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__1__21_chanx_left_out[0:29]),
		.ccff_tail(sb_1__1__21_ccff_tail));

	sb_1__1_ sb_4__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__26_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__29_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__25_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_25_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__22_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_25_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_18_ccff_tail),
		.chany_top_out(sb_1__1__22_chany_top_out[0:29]),
		.chanx_right_out(sb_1__1__22_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__1__22_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__1__22_chanx_left_out[0:29]),
		.ccff_tail(sb_1__1__22_ccff_tail));

	sb_1__1_ sb_4__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__27_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__30_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__26_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_26_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__23_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_26_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_35_ccff_tail),
		.chany_top_out(sb_1__1__23_chany_top_out[0:29]),
		.chanx_right_out(sb_1__1__23_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__1__23_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__1__23_chanx_left_out[0:29]),
		.ccff_tail(sb_1__1__23_ccff_tail));

	sb_1__1_ sb_4__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__28_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__31_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__27_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_27_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__24_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_27_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_20_ccff_tail),
		.chany_top_out(sb_1__1__24_chany_top_out[0:29]),
		.chanx_right_out(sb_1__1__24_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__1__24_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__1__24_chanx_left_out[0:29]),
		.ccff_tail(sb_1__1__24_ccff_tail));

	sb_1__1_ sb_4__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__29_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__32_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__28_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_28_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__25_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_28_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_37_ccff_tail),
		.chany_top_out(sb_1__1__25_chany_top_out[0:29]),
		.chanx_right_out(sb_1__1__25_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__1__25_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__1__25_chanx_left_out[0:29]),
		.ccff_tail(sb_1__1__25_ccff_tail));

	sb_1__1_ sb_4__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__30_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__33_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__29_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_29_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__26_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_29_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_22_ccff_tail),
		.chany_top_out(sb_1__1__26_chany_top_out[0:29]),
		.chanx_right_out(sb_1__1__26_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__1__26_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__1__26_chanx_left_out[0:29]),
		.ccff_tail(sb_1__1__26_ccff_tail));

	sb_1__1_ sb_4__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__31_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__34_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__30_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_30_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__27_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_30_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_39_ccff_tail),
		.chany_top_out(sb_1__1__27_chany_top_out[0:29]),
		.chanx_right_out(sb_1__1__27_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__1__27_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__1__27_chanx_left_out[0:29]),
		.ccff_tail(sb_1__1__27_ccff_tail));

	sb_1__1_ sb_5__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__33_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__35_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__32_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_32_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__28_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_32_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_41_ccff_tail),
		.chany_top_out(sb_1__1__28_chany_top_out[0:29]),
		.chanx_right_out(sb_1__1__28_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__1__28_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__1__28_chanx_left_out[0:29]),
		.ccff_tail(sb_1__1__28_ccff_tail));

	sb_1__1_ sb_5__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__34_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__36_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__33_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_33_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__29_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_33_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_26_ccff_tail),
		.chany_top_out(sb_1__1__29_chany_top_out[0:29]),
		.chanx_right_out(sb_1__1__29_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__1__29_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__1__29_chanx_left_out[0:29]),
		.ccff_tail(sb_1__1__29_ccff_tail));

	sb_1__1_ sb_5__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__35_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__37_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__34_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_34_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__30_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_34_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_43_ccff_tail),
		.chany_top_out(sb_1__1__30_chany_top_out[0:29]),
		.chanx_right_out(sb_1__1__30_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__1__30_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__1__30_chanx_left_out[0:29]),
		.ccff_tail(sb_1__1__30_ccff_tail));

	sb_1__1_ sb_5__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__36_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__38_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__35_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_35_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__31_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_35_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_28_ccff_tail),
		.chany_top_out(sb_1__1__31_chany_top_out[0:29]),
		.chanx_right_out(sb_1__1__31_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__1__31_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__1__31_chanx_left_out[0:29]),
		.ccff_tail(sb_1__1__31_ccff_tail));

	sb_1__1_ sb_5__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__37_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__39_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__36_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_36_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__32_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_36_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_45_ccff_tail),
		.chany_top_out(sb_1__1__32_chany_top_out[0:29]),
		.chanx_right_out(sb_1__1__32_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__1__32_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__1__32_chanx_left_out[0:29]),
		.ccff_tail(sb_1__1__32_ccff_tail));

	sb_1__1_ sb_5__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__38_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__40_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__37_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_37_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__33_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_37_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_30_ccff_tail),
		.chany_top_out(sb_1__1__33_chany_top_out[0:29]),
		.chanx_right_out(sb_1__1__33_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__1__33_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__1__33_chanx_left_out[0:29]),
		.ccff_tail(sb_1__1__33_ccff_tail));

	sb_1__1_ sb_5__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__39_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__41_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__38_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_38_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__34_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_38_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_47_ccff_tail),
		.chany_top_out(sb_1__1__34_chany_top_out[0:29]),
		.chanx_right_out(sb_1__1__34_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__1__34_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__1__34_chanx_left_out[0:29]),
		.ccff_tail(sb_1__1__34_ccff_tail));

	sb_1__1_ sb_6__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__41_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__42_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__40_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_40_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__35_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_40_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_49_ccff_tail),
		.chany_top_out(sb_1__1__35_chany_top_out[0:29]),
		.chanx_right_out(sb_1__1__35_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__1__35_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__1__35_chanx_left_out[0:29]),
		.ccff_tail(sb_1__1__35_ccff_tail));

	sb_1__1_ sb_6__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__42_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__43_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__41_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_41_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__36_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_41_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_34_ccff_tail),
		.chany_top_out(sb_1__1__36_chany_top_out[0:29]),
		.chanx_right_out(sb_1__1__36_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__1__36_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__1__36_chanx_left_out[0:29]),
		.ccff_tail(sb_1__1__36_ccff_tail));

	sb_1__1_ sb_6__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__43_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__44_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__42_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_42_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__37_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_42_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_51_ccff_tail),
		.chany_top_out(sb_1__1__37_chany_top_out[0:29]),
		.chanx_right_out(sb_1__1__37_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__1__37_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__1__37_chanx_left_out[0:29]),
		.ccff_tail(sb_1__1__37_ccff_tail));

	sb_1__1_ sb_6__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__44_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__45_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__43_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_43_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__38_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_43_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_36_ccff_tail),
		.chany_top_out(sb_1__1__38_chany_top_out[0:29]),
		.chanx_right_out(sb_1__1__38_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__1__38_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__1__38_chanx_left_out[0:29]),
		.ccff_tail(sb_1__1__38_ccff_tail));

	sb_1__1_ sb_6__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__45_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__46_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__44_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_44_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__39_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_44_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_53_ccff_tail),
		.chany_top_out(sb_1__1__39_chany_top_out[0:29]),
		.chanx_right_out(sb_1__1__39_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__1__39_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__1__39_chanx_left_out[0:29]),
		.ccff_tail(sb_1__1__39_ccff_tail));

	sb_1__1_ sb_6__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__46_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__47_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__45_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_45_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__40_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_45_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_38_ccff_tail),
		.chany_top_out(sb_1__1__40_chany_top_out[0:29]),
		.chanx_right_out(sb_1__1__40_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__1__40_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__1__40_chanx_left_out[0:29]),
		.ccff_tail(sb_1__1__40_ccff_tail));

	sb_1__1_ sb_6__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__47_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__48_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__46_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_46_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__41_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_46_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_55_ccff_tail),
		.chany_top_out(sb_1__1__41_chany_top_out[0:29]),
		.chanx_right_out(sb_1__1__41_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__1__41_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__1__41_chanx_left_out[0:29]),
		.ccff_tail(sb_1__1__41_ccff_tail));

	sb_1__1_ sb_7__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__49_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__49_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__48_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_48_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__42_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_48_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_57_ccff_tail),
		.chany_top_out(sb_1__1__42_chany_top_out[0:29]),
		.chanx_right_out(sb_1__1__42_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__1__42_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__1__42_chanx_left_out[0:29]),
		.ccff_tail(sb_1__1__42_ccff_tail));

	sb_1__1_ sb_7__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__50_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__50_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__49_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_49_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__43_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_49_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_42_ccff_tail),
		.chany_top_out(sb_1__1__43_chany_top_out[0:29]),
		.chanx_right_out(sb_1__1__43_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__1__43_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__1__43_chanx_left_out[0:29]),
		.ccff_tail(sb_1__1__43_ccff_tail));

	sb_1__1_ sb_7__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__51_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__51_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__50_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_50_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__44_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_50_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_59_ccff_tail),
		.chany_top_out(sb_1__1__44_chany_top_out[0:29]),
		.chanx_right_out(sb_1__1__44_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__1__44_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__1__44_chanx_left_out[0:29]),
		.ccff_tail(sb_1__1__44_ccff_tail));

	sb_1__1_ sb_7__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__52_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__52_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__51_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_51_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__45_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_51_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_44_ccff_tail),
		.chany_top_out(sb_1__1__45_chany_top_out[0:29]),
		.chanx_right_out(sb_1__1__45_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__1__45_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__1__45_chanx_left_out[0:29]),
		.ccff_tail(sb_1__1__45_ccff_tail));

	sb_1__1_ sb_7__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__53_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__53_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__52_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_52_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__46_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_52_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_61_ccff_tail),
		.chany_top_out(sb_1__1__46_chany_top_out[0:29]),
		.chanx_right_out(sb_1__1__46_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__1__46_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__1__46_chanx_left_out[0:29]),
		.ccff_tail(sb_1__1__46_ccff_tail));

	sb_1__1_ sb_7__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__54_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__54_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__53_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_53_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__47_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_53_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_46_ccff_tail),
		.chany_top_out(sb_1__1__47_chany_top_out[0:29]),
		.chanx_right_out(sb_1__1__47_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__1__47_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__1__47_chanx_left_out[0:29]),
		.ccff_tail(sb_1__1__47_ccff_tail));

	sb_1__1_ sb_7__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_1__1__55_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_right_in(cbx_1__1__55_chanx_left_out[0:29]),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__54_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_54_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__48_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_54_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_63_ccff_tail),
		.chany_top_out(sb_1__1__48_chany_top_out[0:29]),
		.chanx_right_out(sb_1__1__48_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__1__48_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__1__48_chanx_left_out[0:29]),
		.ccff_tail(sb_1__1__48_ccff_tail));

	sb_1__8_ sb_1__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__8__1_chanx_left_out[0:29]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_top_1_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_top_1_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_top_1_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__7_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_7_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__8__0_chanx_right_out[0:29]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_0_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_top_0_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_top_0_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_top_0_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_7_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_io_top_top_1_ccff_tail),
		.chanx_right_out(sb_1__8__0_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__8__0_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__8__0_chanx_left_out[0:29]),
		.ccff_tail(sb_1__8__0_ccff_tail));

	sb_1__8_ sb_2__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__8__2_chanx_left_out[0:29]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_top_2_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_top_2_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_top_2_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__15_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_15_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__8__1_chanx_right_out[0:29]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_1_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_top_1_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_top_1_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_top_1_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_15_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_io_top_top_2_ccff_tail),
		.chanx_right_out(sb_1__8__1_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__8__1_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__8__1_chanx_left_out[0:29]),
		.ccff_tail(sb_1__8__1_ccff_tail));

	sb_1__8_ sb_3__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__8__3_chanx_left_out[0:29]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_top_3_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_top_3_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_top_3_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__23_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_23_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__8__2_chanx_right_out[0:29]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_2_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_top_2_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_top_2_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_top_2_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_23_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_io_top_top_3_ccff_tail),
		.chanx_right_out(sb_1__8__2_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__8__2_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__8__2_chanx_left_out[0:29]),
		.ccff_tail(sb_1__8__2_ccff_tail));

	sb_1__8_ sb_4__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__8__4_chanx_left_out[0:29]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_4_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_top_4_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_top_4_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_top_4_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__31_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_31_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__8__3_chanx_right_out[0:29]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_3_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_top_3_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_top_3_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_top_3_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_31_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_io_top_top_4_ccff_tail),
		.chanx_right_out(sb_1__8__3_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__8__3_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__8__3_chanx_left_out[0:29]),
		.ccff_tail(sb_1__8__3_ccff_tail));

	sb_1__8_ sb_5__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__8__5_chanx_left_out[0:29]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_5_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_top_5_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_top_5_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_top_5_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__39_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_39_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__8__4_chanx_right_out[0:29]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_4_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_top_4_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_top_4_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_top_4_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_39_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_io_top_top_5_ccff_tail),
		.chanx_right_out(sb_1__8__4_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__8__4_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__8__4_chanx_left_out[0:29]),
		.ccff_tail(sb_1__8__4_ccff_tail));

	sb_1__8_ sb_6__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__8__6_chanx_left_out[0:29]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_6_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_top_6_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_top_6_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_top_6_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__47_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_47_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__8__5_chanx_right_out[0:29]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_5_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_top_5_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_top_5_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_top_5_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_47_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_io_top_top_6_ccff_tail),
		.chanx_right_out(sb_1__8__5_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__8__5_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__8__5_chanx_left_out[0:29]),
		.ccff_tail(sb_1__8__5_ccff_tail));

	sb_1__8_ sb_7__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_right_in(cbx_1__8__7_chanx_left_out[0:29]),
		.right_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_7_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_top_7_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_top_7_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.right_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_top_7_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_0_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_1_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_2_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_3_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_4_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_5_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_6_),
		.right_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_7_),
		.chany_bottom_in(cby_1__1__55_chany_top_out[0:29]),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_55_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__8__6_chanx_right_out[0:29]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_6_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_top_6_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_top_6_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_top_6_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_55_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_io_top_top_7_ccff_tail),
		.chanx_right_out(sb_1__8__6_chanx_right_out[0:29]),
		.chany_bottom_out(sb_1__8__6_chany_bottom_out[0:29]),
		.chanx_left_out(sb_1__8__6_chanx_left_out[0:29]),
		.ccff_tail(sb_1__8__6_ccff_tail));

	sb_8__0_ sb_8__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_8__1__0_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_7_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_right_7_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_right_7_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_right_7_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.chanx_left_in(cbx_1__0__7_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_bottom_bottom_0_top_width_0_height_0_subtile_3__pin_inpad_0_),
		.ccff_head(grid_clb_48_ccff_tail),
		.chany_top_out(sb_8__0__0_chany_top_out[0:29]),
		.chanx_left_out(sb_8__0__0_chanx_left_out[0:29]),
		.ccff_tail(sb_8__0__0_ccff_tail));

	sb_8__1_ sb_8__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_8__1__1_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_6_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_right_6_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_right_6_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_right_6_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.chany_bottom_in(cby_8__1__0_chany_top_out[0:29]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_7_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_right_7_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_right_7_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_right_7_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_56_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__49_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_56_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_56_ccff_tail),
		.chany_top_out(sb_8__1__0_chany_top_out[0:29]),
		.chany_bottom_out(sb_8__1__0_chany_bottom_out[0:29]),
		.chanx_left_out(sb_8__1__0_chanx_left_out[0:29]),
		.ccff_tail(sb_8__1__0_ccff_tail));

	sb_8__1_ sb_8__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_8__1__2_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_5_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_right_5_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_right_5_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_right_5_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.chany_bottom_in(cby_8__1__1_chany_top_out[0:29]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_6_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_right_6_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_right_6_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_right_6_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_57_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__50_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_57_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_50_ccff_tail),
		.chany_top_out(sb_8__1__1_chany_top_out[0:29]),
		.chany_bottom_out(sb_8__1__1_chany_bottom_out[0:29]),
		.chanx_left_out(sb_8__1__1_chanx_left_out[0:29]),
		.ccff_tail(sb_8__1__1_ccff_tail));

	sb_8__1_ sb_8__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_8__1__3_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_4_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_right_4_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_right_4_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_right_4_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.chany_bottom_in(cby_8__1__2_chany_top_out[0:29]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_5_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_right_5_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_right_5_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_right_5_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_58_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__51_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_58_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_58_ccff_tail),
		.chany_top_out(sb_8__1__2_chany_top_out[0:29]),
		.chany_bottom_out(sb_8__1__2_chany_bottom_out[0:29]),
		.chanx_left_out(sb_8__1__2_chanx_left_out[0:29]),
		.ccff_tail(sb_8__1__2_ccff_tail));

	sb_8__1_ sb_8__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_8__1__4_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_3_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_right_3_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_right_3_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_right_3_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.chany_bottom_in(cby_8__1__3_chany_top_out[0:29]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_4_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_right_4_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_right_4_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_right_4_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_59_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__52_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_59_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_52_ccff_tail),
		.chany_top_out(sb_8__1__3_chany_top_out[0:29]),
		.chany_bottom_out(sb_8__1__3_chany_bottom_out[0:29]),
		.chanx_left_out(sb_8__1__3_chanx_left_out[0:29]),
		.ccff_tail(sb_8__1__3_ccff_tail));

	sb_8__1_ sb_8__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_8__1__5_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_right_2_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_right_2_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_right_2_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.chany_bottom_in(cby_8__1__4_chany_top_out[0:29]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_3_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_right_3_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_right_3_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_right_3_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_60_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__53_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_60_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_60_ccff_tail),
		.chany_top_out(sb_8__1__4_chany_top_out[0:29]),
		.chany_bottom_out(sb_8__1__4_chany_bottom_out[0:29]),
		.chanx_left_out(sb_8__1__4_chanx_left_out[0:29]),
		.ccff_tail(sb_8__1__4_ccff_tail));

	sb_8__1_ sb_8__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_8__1__6_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_right_1_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_right_1_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_right_1_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.chany_bottom_in(cby_8__1__5_chany_top_out[0:29]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_2_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_right_2_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_right_2_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_right_2_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_61_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__54_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_61_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_54_ccff_tail),
		.chany_top_out(sb_8__1__5_chany_top_out[0:29]),
		.chany_bottom_out(sb_8__1__5_chany_bottom_out[0:29]),
		.chanx_left_out(sb_8__1__5_chanx_left_out[0:29]),
		.ccff_tail(sb_8__1__5_ccff_tail));

	sb_8__1_ sb_8__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_top_in(cby_8__1__7_chany_bottom_out[0:29]),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_8_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_9_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_10_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_11_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_12_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_13_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_14_),
		.top_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_15_),
		.top_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_right_0_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_right_0_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.top_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_right_0_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.chany_bottom_in(cby_8__1__6_chany_top_out[0:29]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_1_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_right_1_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_right_1_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_right_1_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_62_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__1__55_chanx_right_out[0:29]),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_62_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_clb_62_ccff_tail),
		.chany_top_out(sb_8__1__6_chany_top_out[0:29]),
		.chany_bottom_out(sb_8__1__6_chany_bottom_out[0:29]),
		.chanx_left_out(sb_8__1__6_chanx_left_out[0:29]),
		.ccff_tail(sb_8__1__6_ccff_tail));

	sb_8__8_ sb_8__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(cby_8__1__7_chany_top_out[0:29]),
		.bottom_right_grid_left_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_right_right_0_left_width_0_height_0_subtile_0__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_right_right_0_left_width_0_height_0_subtile_1__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_right_right_0_left_width_0_height_0_subtile_2__pin_inpad_0_),
		.bottom_right_grid_left_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_right_right_0_left_width_0_height_0_subtile_3__pin_inpad_0_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_8_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_8_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_9_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_9_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_10_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_10_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_11_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_11_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_12_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_12_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_13_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_13_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_14_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_14_),
		.bottom_left_grid_right_width_0_height_0_subtile_0__pin_O_15_(grid_clb_63_right_width_0_height_0_subtile_0__pin_O_15_),
		.chanx_left_in(cbx_1__8__7_chanx_right_out[0:29]),
		.left_top_grid_bottom_width_0_height_0_subtile_0__pin_inpad_0_(grid_io_top_top_7_bottom_width_0_height_0_subtile_0__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_1__pin_inpad_0_(grid_io_top_top_7_bottom_width_0_height_0_subtile_1__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_2__pin_inpad_0_(grid_io_top_top_7_bottom_width_0_height_0_subtile_2__pin_inpad_0_),
		.left_top_grid_bottom_width_0_height_0_subtile_3__pin_inpad_0_(grid_io_top_top_7_bottom_width_0_height_0_subtile_3__pin_inpad_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_0_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_0_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_1_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_1_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_2_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_2_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_3_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_3_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_4_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_4_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_5_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_5_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_6_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_6_),
		.left_bottom_grid_top_width_0_height_0_subtile_0__pin_O_7_(grid_clb_63_top_width_0_height_0_subtile_0__pin_O_7_),
		.ccff_head(grid_io_right_right_0_ccff_tail),
		.chany_bottom_out(sb_8__8__0_chany_bottom_out[0:29]),
		.chanx_left_out(sb_8__8__0_chanx_left_out[0:29]),
		.ccff_tail(sb_8__8__0_ccff_tail));

	cbx_1__0_ cbx_1__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__0__0_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__0__0_chanx_left_out[0:29]),
		.ccff_head(sb_1__0__0_ccff_tail),
		.chanx_left_out(cbx_1__0__0_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__0__0_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__0_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.ccff_tail(cbx_1__0__0_ccff_tail));

	cbx_1__0_ cbx_2__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__0_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__0__1_chanx_left_out[0:29]),
		.ccff_head(sb_1__0__1_ccff_tail),
		.chanx_left_out(cbx_1__0__1_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__0__1_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__1_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.ccff_tail(cbx_1__0__1_ccff_tail));

	cbx_1__0_ cbx_3__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__1_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__0__2_chanx_left_out[0:29]),
		.ccff_head(sb_1__0__2_ccff_tail),
		.chanx_left_out(cbx_1__0__2_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__0__2_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__2_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.ccff_tail(cbx_1__0__2_ccff_tail));

	cbx_1__0_ cbx_4__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__2_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__0__3_chanx_left_out[0:29]),
		.ccff_head(sb_1__0__3_ccff_tail),
		.chanx_left_out(cbx_1__0__3_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__0__3_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__3_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.ccff_tail(cbx_1__0__3_ccff_tail));

	cbx_1__0_ cbx_5__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__3_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__0__4_chanx_left_out[0:29]),
		.ccff_head(sb_1__0__4_ccff_tail),
		.chanx_left_out(cbx_1__0__4_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__0__4_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__4_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.ccff_tail(cbx_1__0__4_ccff_tail));

	cbx_1__0_ cbx_6__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__4_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__0__5_chanx_left_out[0:29]),
		.ccff_head(sb_1__0__5_ccff_tail),
		.chanx_left_out(cbx_1__0__5_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__0__5_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__5_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.ccff_tail(cbx_1__0__5_ccff_tail));

	cbx_1__0_ cbx_7__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__5_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__0__6_chanx_left_out[0:29]),
		.ccff_head(sb_1__0__6_ccff_tail),
		.chanx_left_out(cbx_1__0__6_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__0__6_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__6_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.ccff_tail(cbx_1__0__6_ccff_tail));

	cbx_1__0_ cbx_8__0_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__0__6_chanx_right_out[0:29]),
		.chanx_right_in(sb_8__0__0_chanx_left_out[0:29]),
		.ccff_head(sb_8__0__0_ccff_tail),
		.chanx_left_out(cbx_1__0__7_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__0__7_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_0__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_1__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_2__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__0__7_bottom_grid_top_width_0_height_0_subtile_3__pin_outpad_0_),
		.ccff_tail(cbx_1__0__7_ccff_tail));

	cbx_1__1_ cbx_1__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__1__0_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__1__0_chanx_left_out[0:29]),
		.ccff_head(sb_1__1__0_ccff_tail),
		.chanx_left_out(cbx_1__1__0_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__0_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__0_ccff_tail));

	cbx_1__1_ cbx_1__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__1__1_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__1__1_chanx_left_out[0:29]),
		.ccff_head(sb_1__1__1_ccff_tail),
		.chanx_left_out(cbx_1__1__1_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__1_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__1_ccff_tail));

	cbx_1__1_ cbx_1__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__1__2_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__1__2_chanx_left_out[0:29]),
		.ccff_head(sb_1__1__2_ccff_tail),
		.chanx_left_out(cbx_1__1__2_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__2_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__2_ccff_tail));

	cbx_1__1_ cbx_1__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__1__3_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__1__3_chanx_left_out[0:29]),
		.ccff_head(sb_1__1__3_ccff_tail),
		.chanx_left_out(cbx_1__1__3_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__3_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__3_ccff_tail));

	cbx_1__1_ cbx_1__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__1__4_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__1__4_chanx_left_out[0:29]),
		.ccff_head(sb_1__1__4_ccff_tail),
		.chanx_left_out(cbx_1__1__4_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__4_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__4_ccff_tail));

	cbx_1__1_ cbx_1__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__1__5_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__1__5_chanx_left_out[0:29]),
		.ccff_head(sb_1__1__5_ccff_tail),
		.chanx_left_out(cbx_1__1__5_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__5_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__5_ccff_tail));

	cbx_1__1_ cbx_1__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__1__6_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__1__6_chanx_left_out[0:29]),
		.ccff_head(sb_1__1__6_ccff_tail),
		.chanx_left_out(cbx_1__1__6_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__6_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__6_ccff_tail));

	cbx_1__1_ cbx_2__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__0_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__1__7_chanx_left_out[0:29]),
		.ccff_head(sb_1__1__7_ccff_tail),
		.chanx_left_out(cbx_1__1__7_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__7_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__7_ccff_tail));

	cbx_1__1_ cbx_2__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__1_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__1__8_chanx_left_out[0:29]),
		.ccff_head(sb_1__1__8_ccff_tail),
		.chanx_left_out(cbx_1__1__8_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__8_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__8_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__8_ccff_tail));

	cbx_1__1_ cbx_2__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__2_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__1__9_chanx_left_out[0:29]),
		.ccff_head(sb_1__1__9_ccff_tail),
		.chanx_left_out(cbx_1__1__9_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__9_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__9_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__9_ccff_tail));

	cbx_1__1_ cbx_2__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__3_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__1__10_chanx_left_out[0:29]),
		.ccff_head(sb_1__1__10_ccff_tail),
		.chanx_left_out(cbx_1__1__10_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__10_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__10_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__10_ccff_tail));

	cbx_1__1_ cbx_2__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__4_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__1__11_chanx_left_out[0:29]),
		.ccff_head(sb_1__1__11_ccff_tail),
		.chanx_left_out(cbx_1__1__11_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__11_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__11_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__11_ccff_tail));

	cbx_1__1_ cbx_2__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__5_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__1__12_chanx_left_out[0:29]),
		.ccff_head(sb_1__1__12_ccff_tail),
		.chanx_left_out(cbx_1__1__12_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__12_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__12_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__12_ccff_tail));

	cbx_1__1_ cbx_2__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__6_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__1__13_chanx_left_out[0:29]),
		.ccff_head(sb_1__1__13_ccff_tail),
		.chanx_left_out(cbx_1__1__13_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__13_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__13_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__13_ccff_tail));

	cbx_1__1_ cbx_3__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__7_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__1__14_chanx_left_out[0:29]),
		.ccff_head(sb_1__1__14_ccff_tail),
		.chanx_left_out(cbx_1__1__14_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__14_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__14_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__14_ccff_tail));

	cbx_1__1_ cbx_3__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__8_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__1__15_chanx_left_out[0:29]),
		.ccff_head(sb_1__1__15_ccff_tail),
		.chanx_left_out(cbx_1__1__15_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__15_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__15_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__15_ccff_tail));

	cbx_1__1_ cbx_3__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__9_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__1__16_chanx_left_out[0:29]),
		.ccff_head(sb_1__1__16_ccff_tail),
		.chanx_left_out(cbx_1__1__16_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__16_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__16_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__16_ccff_tail));

	cbx_1__1_ cbx_3__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__10_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__1__17_chanx_left_out[0:29]),
		.ccff_head(sb_1__1__17_ccff_tail),
		.chanx_left_out(cbx_1__1__17_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__17_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__17_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__17_ccff_tail));

	cbx_1__1_ cbx_3__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__11_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__1__18_chanx_left_out[0:29]),
		.ccff_head(sb_1__1__18_ccff_tail),
		.chanx_left_out(cbx_1__1__18_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__18_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__18_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__18_ccff_tail));

	cbx_1__1_ cbx_3__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__12_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__1__19_chanx_left_out[0:29]),
		.ccff_head(sb_1__1__19_ccff_tail),
		.chanx_left_out(cbx_1__1__19_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__19_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__19_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__19_ccff_tail));

	cbx_1__1_ cbx_3__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__13_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__1__20_chanx_left_out[0:29]),
		.ccff_head(sb_1__1__20_ccff_tail),
		.chanx_left_out(cbx_1__1__20_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__20_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__20_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__20_ccff_tail));

	cbx_1__1_ cbx_4__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__14_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__1__21_chanx_left_out[0:29]),
		.ccff_head(sb_1__1__21_ccff_tail),
		.chanx_left_out(cbx_1__1__21_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__21_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__21_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__21_ccff_tail));

	cbx_1__1_ cbx_4__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__15_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__1__22_chanx_left_out[0:29]),
		.ccff_head(sb_1__1__22_ccff_tail),
		.chanx_left_out(cbx_1__1__22_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__22_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__22_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__22_ccff_tail));

	cbx_1__1_ cbx_4__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__16_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__1__23_chanx_left_out[0:29]),
		.ccff_head(sb_1__1__23_ccff_tail),
		.chanx_left_out(cbx_1__1__23_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__23_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__23_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__23_ccff_tail));

	cbx_1__1_ cbx_4__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__17_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__1__24_chanx_left_out[0:29]),
		.ccff_head(sb_1__1__24_ccff_tail),
		.chanx_left_out(cbx_1__1__24_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__24_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__24_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__24_ccff_tail));

	cbx_1__1_ cbx_4__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__18_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__1__25_chanx_left_out[0:29]),
		.ccff_head(sb_1__1__25_ccff_tail),
		.chanx_left_out(cbx_1__1__25_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__25_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__25_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__25_ccff_tail));

	cbx_1__1_ cbx_4__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__19_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__1__26_chanx_left_out[0:29]),
		.ccff_head(sb_1__1__26_ccff_tail),
		.chanx_left_out(cbx_1__1__26_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__26_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__26_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__26_ccff_tail));

	cbx_1__1_ cbx_4__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__20_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__1__27_chanx_left_out[0:29]),
		.ccff_head(sb_1__1__27_ccff_tail),
		.chanx_left_out(cbx_1__1__27_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__27_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__27_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__27_ccff_tail));

	cbx_1__1_ cbx_5__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__21_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__1__28_chanx_left_out[0:29]),
		.ccff_head(sb_1__1__28_ccff_tail),
		.chanx_left_out(cbx_1__1__28_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__28_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__28_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__28_ccff_tail));

	cbx_1__1_ cbx_5__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__22_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__1__29_chanx_left_out[0:29]),
		.ccff_head(sb_1__1__29_ccff_tail),
		.chanx_left_out(cbx_1__1__29_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__29_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__29_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__29_ccff_tail));

	cbx_1__1_ cbx_5__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__23_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__1__30_chanx_left_out[0:29]),
		.ccff_head(sb_1__1__30_ccff_tail),
		.chanx_left_out(cbx_1__1__30_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__30_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__30_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__30_ccff_tail));

	cbx_1__1_ cbx_5__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__24_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__1__31_chanx_left_out[0:29]),
		.ccff_head(sb_1__1__31_ccff_tail),
		.chanx_left_out(cbx_1__1__31_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__31_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__31_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__31_ccff_tail));

	cbx_1__1_ cbx_5__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__25_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__1__32_chanx_left_out[0:29]),
		.ccff_head(sb_1__1__32_ccff_tail),
		.chanx_left_out(cbx_1__1__32_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__32_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__32_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__32_ccff_tail));

	cbx_1__1_ cbx_5__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__26_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__1__33_chanx_left_out[0:29]),
		.ccff_head(sb_1__1__33_ccff_tail),
		.chanx_left_out(cbx_1__1__33_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__33_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__33_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__33_ccff_tail));

	cbx_1__1_ cbx_5__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__27_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__1__34_chanx_left_out[0:29]),
		.ccff_head(sb_1__1__34_ccff_tail),
		.chanx_left_out(cbx_1__1__34_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__34_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__34_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__34_ccff_tail));

	cbx_1__1_ cbx_6__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__28_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__1__35_chanx_left_out[0:29]),
		.ccff_head(sb_1__1__35_ccff_tail),
		.chanx_left_out(cbx_1__1__35_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__35_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__35_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__35_ccff_tail));

	cbx_1__1_ cbx_6__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__29_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__1__36_chanx_left_out[0:29]),
		.ccff_head(sb_1__1__36_ccff_tail),
		.chanx_left_out(cbx_1__1__36_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__36_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__36_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__36_ccff_tail));

	cbx_1__1_ cbx_6__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__30_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__1__37_chanx_left_out[0:29]),
		.ccff_head(sb_1__1__37_ccff_tail),
		.chanx_left_out(cbx_1__1__37_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__37_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__37_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__37_ccff_tail));

	cbx_1__1_ cbx_6__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__31_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__1__38_chanx_left_out[0:29]),
		.ccff_head(sb_1__1__38_ccff_tail),
		.chanx_left_out(cbx_1__1__38_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__38_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__38_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__38_ccff_tail));

	cbx_1__1_ cbx_6__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__32_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__1__39_chanx_left_out[0:29]),
		.ccff_head(sb_1__1__39_ccff_tail),
		.chanx_left_out(cbx_1__1__39_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__39_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__39_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__39_ccff_tail));

	cbx_1__1_ cbx_6__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__33_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__1__40_chanx_left_out[0:29]),
		.ccff_head(sb_1__1__40_ccff_tail),
		.chanx_left_out(cbx_1__1__40_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__40_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__40_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__40_ccff_tail));

	cbx_1__1_ cbx_6__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__34_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__1__41_chanx_left_out[0:29]),
		.ccff_head(sb_1__1__41_ccff_tail),
		.chanx_left_out(cbx_1__1__41_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__41_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__41_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__41_ccff_tail));

	cbx_1__1_ cbx_7__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__35_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__1__42_chanx_left_out[0:29]),
		.ccff_head(sb_1__1__42_ccff_tail),
		.chanx_left_out(cbx_1__1__42_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__42_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__42_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__42_ccff_tail));

	cbx_1__1_ cbx_7__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__36_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__1__43_chanx_left_out[0:29]),
		.ccff_head(sb_1__1__43_ccff_tail),
		.chanx_left_out(cbx_1__1__43_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__43_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__43_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__43_ccff_tail));

	cbx_1__1_ cbx_7__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__37_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__1__44_chanx_left_out[0:29]),
		.ccff_head(sb_1__1__44_ccff_tail),
		.chanx_left_out(cbx_1__1__44_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__44_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__44_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__44_ccff_tail));

	cbx_1__1_ cbx_7__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__38_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__1__45_chanx_left_out[0:29]),
		.ccff_head(sb_1__1__45_ccff_tail),
		.chanx_left_out(cbx_1__1__45_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__45_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__45_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__45_ccff_tail));

	cbx_1__1_ cbx_7__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__39_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__1__46_chanx_left_out[0:29]),
		.ccff_head(sb_1__1__46_ccff_tail),
		.chanx_left_out(cbx_1__1__46_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__46_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__46_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__46_ccff_tail));

	cbx_1__1_ cbx_7__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__40_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__1__47_chanx_left_out[0:29]),
		.ccff_head(sb_1__1__47_ccff_tail),
		.chanx_left_out(cbx_1__1__47_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__47_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__47_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__47_ccff_tail));

	cbx_1__1_ cbx_7__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__41_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__1__48_chanx_left_out[0:29]),
		.ccff_head(sb_1__1__48_ccff_tail),
		.chanx_left_out(cbx_1__1__48_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__48_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__48_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__48_ccff_tail));

	cbx_1__1_ cbx_8__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__42_chanx_right_out[0:29]),
		.chanx_right_in(sb_8__1__0_chanx_left_out[0:29]),
		.ccff_head(sb_8__1__0_ccff_tail),
		.chanx_left_out(cbx_1__1__49_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__49_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__49_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__49_ccff_tail));

	cbx_1__1_ cbx_8__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__43_chanx_right_out[0:29]),
		.chanx_right_in(sb_8__1__1_chanx_left_out[0:29]),
		.ccff_head(sb_8__1__1_ccff_tail),
		.chanx_left_out(cbx_1__1__50_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__50_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__50_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__50_ccff_tail));

	cbx_1__1_ cbx_8__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__44_chanx_right_out[0:29]),
		.chanx_right_in(sb_8__1__2_chanx_left_out[0:29]),
		.ccff_head(sb_8__1__2_ccff_tail),
		.chanx_left_out(cbx_1__1__51_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__51_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__51_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__51_ccff_tail));

	cbx_1__1_ cbx_8__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__45_chanx_right_out[0:29]),
		.chanx_right_in(sb_8__1__3_chanx_left_out[0:29]),
		.ccff_head(sb_8__1__3_ccff_tail),
		.chanx_left_out(cbx_1__1__52_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__52_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__52_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__52_ccff_tail));

	cbx_1__1_ cbx_8__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__46_chanx_right_out[0:29]),
		.chanx_right_in(sb_8__1__4_chanx_left_out[0:29]),
		.ccff_head(sb_8__1__4_ccff_tail),
		.chanx_left_out(cbx_1__1__53_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__53_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__53_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__53_ccff_tail));

	cbx_1__1_ cbx_8__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__47_chanx_right_out[0:29]),
		.chanx_right_in(sb_8__1__5_chanx_left_out[0:29]),
		.ccff_head(sb_8__1__5_ccff_tail),
		.chanx_left_out(cbx_1__1__54_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__54_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__54_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__54_ccff_tail));

	cbx_1__1_ cbx_8__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__1__48_chanx_right_out[0:29]),
		.chanx_right_in(sb_8__1__6_chanx_left_out[0:29]),
		.ccff_head(sb_8__1__6_ccff_tail),
		.chanx_left_out(cbx_1__1__55_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__1__55_chanx_right_out[0:29]),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__1__55_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__1__55_ccff_tail));

	cbx_1__8_ cbx_1__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_0__8__0_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__8__0_chanx_left_out[0:29]),
		.ccff_head(sb_1__8__0_ccff_tail),
		.chanx_left_out(cbx_1__8__0_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__8__0_chanx_right_out[0:29]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__8__0_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__8__0_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__8__0_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__8__0_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__8__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__8__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__8__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__8__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__8__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__8__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__8__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__8__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__8__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__8__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__8__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__8__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__8__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__8__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__8__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__8__0_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__8__0_ccff_tail));

	cbx_1__8_ cbx_2__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__8__0_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__8__1_chanx_left_out[0:29]),
		.ccff_head(sb_1__8__1_ccff_tail),
		.chanx_left_out(cbx_1__8__1_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__8__1_chanx_right_out[0:29]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__8__1_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__8__1_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__8__1_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__8__1_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__8__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__8__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__8__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__8__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__8__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__8__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__8__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__8__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__8__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__8__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__8__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__8__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__8__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__8__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__8__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__8__1_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__8__1_ccff_tail));

	cbx_1__8_ cbx_3__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__8__1_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__8__2_chanx_left_out[0:29]),
		.ccff_head(sb_1__8__2_ccff_tail),
		.chanx_left_out(cbx_1__8__2_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__8__2_chanx_right_out[0:29]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__8__2_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__8__2_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__8__2_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__8__2_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__8__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__8__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__8__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__8__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__8__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__8__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__8__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__8__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__8__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__8__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__8__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__8__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__8__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__8__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__8__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__8__2_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__8__2_ccff_tail));

	cbx_1__8_ cbx_4__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__8__2_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__8__3_chanx_left_out[0:29]),
		.ccff_head(sb_1__8__3_ccff_tail),
		.chanx_left_out(cbx_1__8__3_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__8__3_chanx_right_out[0:29]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__8__3_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__8__3_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__8__3_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__8__3_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__8__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__8__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__8__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__8__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__8__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__8__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__8__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__8__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__8__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__8__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__8__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__8__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__8__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__8__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__8__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__8__3_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__8__3_ccff_tail));

	cbx_1__8_ cbx_5__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__8__3_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__8__4_chanx_left_out[0:29]),
		.ccff_head(sb_1__8__4_ccff_tail),
		.chanx_left_out(cbx_1__8__4_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__8__4_chanx_right_out[0:29]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__8__4_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__8__4_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__8__4_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__8__4_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__8__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__8__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__8__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__8__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__8__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__8__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__8__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__8__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__8__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__8__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__8__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__8__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__8__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__8__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__8__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__8__4_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__8__4_ccff_tail));

	cbx_1__8_ cbx_6__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__8__4_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__8__5_chanx_left_out[0:29]),
		.ccff_head(sb_1__8__5_ccff_tail),
		.chanx_left_out(cbx_1__8__5_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__8__5_chanx_right_out[0:29]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__8__5_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__8__5_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__8__5_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__8__5_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__8__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__8__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__8__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__8__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__8__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__8__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__8__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__8__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__8__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__8__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__8__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__8__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__8__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__8__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__8__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__8__5_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__8__5_ccff_tail));

	cbx_1__8_ cbx_7__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__8__5_chanx_right_out[0:29]),
		.chanx_right_in(sb_1__8__6_chanx_left_out[0:29]),
		.ccff_head(sb_1__8__6_ccff_tail),
		.chanx_left_out(cbx_1__8__6_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__8__6_chanx_right_out[0:29]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__8__6_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__8__6_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__8__6_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__8__6_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__8__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__8__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__8__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__8__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__8__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__8__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__8__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__8__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__8__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__8__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__8__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__8__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__8__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__8__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__8__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__8__6_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__8__6_ccff_tail));

	cbx_1__8_ cbx_8__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chanx_left_in(sb_1__8__6_chanx_right_out[0:29]),
		.chanx_right_in(sb_8__8__0_chanx_left_out[0:29]),
		.ccff_head(sb_8__8__0_ccff_tail),
		.chanx_left_out(cbx_1__8__7_chanx_left_out[0:29]),
		.chanx_right_out(cbx_1__8__7_chanx_right_out[0:29]),
		.top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_(cbx_1__8__7_top_grid_bottom_width_0_height_0_subtile_0__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_(cbx_1__8__7_top_grid_bottom_width_0_height_0_subtile_1__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_(cbx_1__8__7_top_grid_bottom_width_0_height_0_subtile_2__pin_outpad_0_),
		.top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_(cbx_1__8__7_top_grid_bottom_width_0_height_0_subtile_3__pin_outpad_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_(cbx_1__8__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_(cbx_1__8__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_(cbx_1__8__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_(cbx_1__8__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I0i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_(cbx_1__8__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_(cbx_1__8__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_(cbx_1__8__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_(cbx_1__8__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I1i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_(cbx_1__8__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_(cbx_1__8__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I2_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_(cbx_1__8__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_(cbx_1__8__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I2i_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_(cbx_1__8__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_(cbx_1__8__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I3_1_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_(cbx_1__8__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_0_),
		.bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_(cbx_1__8__7_bottom_grid_top_width_0_height_0_subtile_0__pin_I3i_1_),
		.ccff_tail(cbx_1__8__7_ccff_tail));

	cby_0__1_ cby_0__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__0__0_chany_top_out[0:29]),
		.chany_top_in(sb_0__1__0_chany_bottom_out[0:29]),
		.ccff_head(sb_0__0__0_ccff_tail),
		.chany_bottom_out(cby_0__1__0_chany_bottom_out[0:29]),
		.chany_top_out(cby_0__1__0_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__0_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.ccff_tail(cby_0__1__0_ccff_tail));

	cby_0__1_ cby_0__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__0_chany_top_out[0:29]),
		.chany_top_in(sb_0__1__1_chany_bottom_out[0:29]),
		.ccff_head(sb_0__1__0_ccff_tail),
		.chany_bottom_out(cby_0__1__1_chany_bottom_out[0:29]),
		.chany_top_out(cby_0__1__1_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__1_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.ccff_tail(cby_0__1__1_ccff_tail));

	cby_0__1_ cby_0__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__1_chany_top_out[0:29]),
		.chany_top_in(sb_0__1__2_chany_bottom_out[0:29]),
		.ccff_head(sb_0__1__1_ccff_tail),
		.chany_bottom_out(cby_0__1__2_chany_bottom_out[0:29]),
		.chany_top_out(cby_0__1__2_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__2_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.ccff_tail(cby_0__1__2_ccff_tail));

	cby_0__1_ cby_0__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__2_chany_top_out[0:29]),
		.chany_top_in(sb_0__1__3_chany_bottom_out[0:29]),
		.ccff_head(sb_0__1__2_ccff_tail),
		.chany_bottom_out(cby_0__1__3_chany_bottom_out[0:29]),
		.chany_top_out(cby_0__1__3_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__3_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.ccff_tail(cby_0__1__3_ccff_tail));

	cby_0__1_ cby_0__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__3_chany_top_out[0:29]),
		.chany_top_in(sb_0__1__4_chany_bottom_out[0:29]),
		.ccff_head(sb_0__1__3_ccff_tail),
		.chany_bottom_out(cby_0__1__4_chany_bottom_out[0:29]),
		.chany_top_out(cby_0__1__4_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__4_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.ccff_tail(cby_0__1__4_ccff_tail));

	cby_0__1_ cby_0__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__4_chany_top_out[0:29]),
		.chany_top_in(sb_0__1__5_chany_bottom_out[0:29]),
		.ccff_head(sb_0__1__4_ccff_tail),
		.chany_bottom_out(cby_0__1__5_chany_bottom_out[0:29]),
		.chany_top_out(cby_0__1__5_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__5_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__5_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__5_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__5_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.ccff_tail(cby_0__1__5_ccff_tail));

	cby_0__1_ cby_0__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__5_chany_top_out[0:29]),
		.chany_top_in(sb_0__1__6_chany_bottom_out[0:29]),
		.ccff_head(sb_0__1__5_ccff_tail),
		.chany_bottom_out(cby_0__1__6_chany_bottom_out[0:29]),
		.chany_top_out(cby_0__1__6_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__6_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__6_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__6_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__6_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.ccff_tail(cby_0__1__6_ccff_tail));

	cby_0__1_ cby_0__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_0__1__6_chany_top_out[0:29]),
		.chany_top_in(sb_0__8__0_chany_bottom_out[0:29]),
		.ccff_head(sb_0__1__6_ccff_tail),
		.chany_bottom_out(cby_0__1__7_chany_bottom_out[0:29]),
		.chany_top_out(cby_0__1__7_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_(cby_0__1__7_left_grid_right_width_0_height_0_subtile_0__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_(cby_0__1__7_left_grid_right_width_0_height_0_subtile_1__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_(cby_0__1__7_left_grid_right_width_0_height_0_subtile_2__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_(cby_0__1__7_left_grid_right_width_0_height_0_subtile_3__pin_outpad_0_),
		.ccff_tail(cby_0__1__7_ccff_tail));

	cby_1__1_ cby_1__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__0__0_chany_top_out[0:29]),
		.chany_top_in(sb_1__1__0_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__0__0_ccff_tail),
		.chany_bottom_out(cby_1__1__0_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__0_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__0_ccff_tail));

	cby_1__1_ cby_1__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__0_chany_top_out[0:29]),
		.chany_top_in(sb_1__1__1_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__0_ccff_tail),
		.chany_bottom_out(cby_1__1__1_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__1_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__1_ccff_tail));

	cby_1__1_ cby_1__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__1_chany_top_out[0:29]),
		.chany_top_in(sb_1__1__2_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__1_ccff_tail),
		.chany_bottom_out(cby_1__1__2_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__2_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__2_ccff_tail));

	cby_1__1_ cby_1__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__2_chany_top_out[0:29]),
		.chany_top_in(sb_1__1__3_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__2_ccff_tail),
		.chany_bottom_out(cby_1__1__3_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__3_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__3_ccff_tail));

	cby_1__1_ cby_1__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__3_chany_top_out[0:29]),
		.chany_top_in(sb_1__1__4_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__3_ccff_tail),
		.chany_bottom_out(cby_1__1__4_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__4_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__4_ccff_tail));

	cby_1__1_ cby_1__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__4_chany_top_out[0:29]),
		.chany_top_in(sb_1__1__5_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__4_ccff_tail),
		.chany_bottom_out(cby_1__1__5_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__5_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__5_ccff_tail));

	cby_1__1_ cby_1__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__5_chany_top_out[0:29]),
		.chany_top_in(sb_1__1__6_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__5_ccff_tail),
		.chany_bottom_out(cby_1__1__6_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__6_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__6_ccff_tail));

	cby_1__1_ cby_1__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__6_chany_top_out[0:29]),
		.chany_top_in(sb_1__8__0_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__6_ccff_tail),
		.chany_bottom_out(cby_1__1__7_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__7_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__7_ccff_tail));

	cby_1__1_ cby_2__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__0__1_chany_top_out[0:29]),
		.chany_top_in(sb_1__1__7_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__0__1_ccff_tail),
		.chany_bottom_out(cby_1__1__8_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__8_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__8_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__8_ccff_tail));

	cby_1__1_ cby_2__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__7_chany_top_out[0:29]),
		.chany_top_in(sb_1__1__8_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__7_ccff_tail),
		.chany_bottom_out(cby_1__1__9_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__9_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__9_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__9_ccff_tail));

	cby_1__1_ cby_2__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__8_chany_top_out[0:29]),
		.chany_top_in(sb_1__1__9_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__8_ccff_tail),
		.chany_bottom_out(cby_1__1__10_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__10_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__10_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__10_ccff_tail));

	cby_1__1_ cby_2__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__9_chany_top_out[0:29]),
		.chany_top_in(sb_1__1__10_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__9_ccff_tail),
		.chany_bottom_out(cby_1__1__11_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__11_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__11_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__11_ccff_tail));

	cby_1__1_ cby_2__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__10_chany_top_out[0:29]),
		.chany_top_in(sb_1__1__11_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__10_ccff_tail),
		.chany_bottom_out(cby_1__1__12_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__12_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__12_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__12_ccff_tail));

	cby_1__1_ cby_2__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__11_chany_top_out[0:29]),
		.chany_top_in(sb_1__1__12_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__11_ccff_tail),
		.chany_bottom_out(cby_1__1__13_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__13_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__13_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__13_ccff_tail));

	cby_1__1_ cby_2__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__12_chany_top_out[0:29]),
		.chany_top_in(sb_1__1__13_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__12_ccff_tail),
		.chany_bottom_out(cby_1__1__14_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__14_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__14_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__14_ccff_tail));

	cby_1__1_ cby_2__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__13_chany_top_out[0:29]),
		.chany_top_in(sb_1__8__1_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__13_ccff_tail),
		.chany_bottom_out(cby_1__1__15_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__15_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__15_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__15_ccff_tail));

	cby_1__1_ cby_3__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__0__2_chany_top_out[0:29]),
		.chany_top_in(sb_1__1__14_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__0__2_ccff_tail),
		.chany_bottom_out(cby_1__1__16_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__16_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__16_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__16_ccff_tail));

	cby_1__1_ cby_3__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__14_chany_top_out[0:29]),
		.chany_top_in(sb_1__1__15_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__14_ccff_tail),
		.chany_bottom_out(cby_1__1__17_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__17_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__17_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__17_ccff_tail));

	cby_1__1_ cby_3__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__15_chany_top_out[0:29]),
		.chany_top_in(sb_1__1__16_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__15_ccff_tail),
		.chany_bottom_out(cby_1__1__18_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__18_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__18_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__18_ccff_tail));

	cby_1__1_ cby_3__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__16_chany_top_out[0:29]),
		.chany_top_in(sb_1__1__17_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__16_ccff_tail),
		.chany_bottom_out(cby_1__1__19_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__19_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__19_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__19_ccff_tail));

	cby_1__1_ cby_3__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__17_chany_top_out[0:29]),
		.chany_top_in(sb_1__1__18_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__17_ccff_tail),
		.chany_bottom_out(cby_1__1__20_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__20_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__20_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__20_ccff_tail));

	cby_1__1_ cby_3__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__18_chany_top_out[0:29]),
		.chany_top_in(sb_1__1__19_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__18_ccff_tail),
		.chany_bottom_out(cby_1__1__21_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__21_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__21_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__21_ccff_tail));

	cby_1__1_ cby_3__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__19_chany_top_out[0:29]),
		.chany_top_in(sb_1__1__20_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__19_ccff_tail),
		.chany_bottom_out(cby_1__1__22_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__22_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__22_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__22_ccff_tail));

	cby_1__1_ cby_3__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__20_chany_top_out[0:29]),
		.chany_top_in(sb_1__8__2_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__20_ccff_tail),
		.chany_bottom_out(cby_1__1__23_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__23_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__23_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__23_ccff_tail));

	cby_1__1_ cby_4__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__0__3_chany_top_out[0:29]),
		.chany_top_in(sb_1__1__21_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__0__3_ccff_tail),
		.chany_bottom_out(cby_1__1__24_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__24_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__24_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__24_ccff_tail));

	cby_1__1_ cby_4__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__21_chany_top_out[0:29]),
		.chany_top_in(sb_1__1__22_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__21_ccff_tail),
		.chany_bottom_out(cby_1__1__25_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__25_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__25_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__25_ccff_tail));

	cby_1__1_ cby_4__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__22_chany_top_out[0:29]),
		.chany_top_in(sb_1__1__23_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__22_ccff_tail),
		.chany_bottom_out(cby_1__1__26_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__26_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__26_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__26_ccff_tail));

	cby_1__1_ cby_4__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__23_chany_top_out[0:29]),
		.chany_top_in(sb_1__1__24_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__23_ccff_tail),
		.chany_bottom_out(cby_1__1__27_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__27_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__27_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__27_ccff_tail));

	cby_1__1_ cby_4__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__24_chany_top_out[0:29]),
		.chany_top_in(sb_1__1__25_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__24_ccff_tail),
		.chany_bottom_out(cby_1__1__28_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__28_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__28_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__28_ccff_tail));

	cby_1__1_ cby_4__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__25_chany_top_out[0:29]),
		.chany_top_in(sb_1__1__26_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__25_ccff_tail),
		.chany_bottom_out(cby_1__1__29_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__29_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__29_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__29_ccff_tail));

	cby_1__1_ cby_4__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__26_chany_top_out[0:29]),
		.chany_top_in(sb_1__1__27_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__26_ccff_tail),
		.chany_bottom_out(cby_1__1__30_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__30_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__30_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__30_ccff_tail));

	cby_1__1_ cby_4__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__27_chany_top_out[0:29]),
		.chany_top_in(sb_1__8__3_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__27_ccff_tail),
		.chany_bottom_out(cby_1__1__31_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__31_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__31_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__31_ccff_tail));

	cby_1__1_ cby_5__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__0__4_chany_top_out[0:29]),
		.chany_top_in(sb_1__1__28_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__0__4_ccff_tail),
		.chany_bottom_out(cby_1__1__32_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__32_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__32_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__32_ccff_tail));

	cby_1__1_ cby_5__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__28_chany_top_out[0:29]),
		.chany_top_in(sb_1__1__29_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__28_ccff_tail),
		.chany_bottom_out(cby_1__1__33_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__33_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__33_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__33_ccff_tail));

	cby_1__1_ cby_5__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__29_chany_top_out[0:29]),
		.chany_top_in(sb_1__1__30_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__29_ccff_tail),
		.chany_bottom_out(cby_1__1__34_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__34_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__34_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__34_ccff_tail));

	cby_1__1_ cby_5__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__30_chany_top_out[0:29]),
		.chany_top_in(sb_1__1__31_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__30_ccff_tail),
		.chany_bottom_out(cby_1__1__35_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__35_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__35_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__35_ccff_tail));

	cby_1__1_ cby_5__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__31_chany_top_out[0:29]),
		.chany_top_in(sb_1__1__32_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__31_ccff_tail),
		.chany_bottom_out(cby_1__1__36_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__36_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__36_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__36_ccff_tail));

	cby_1__1_ cby_5__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__32_chany_top_out[0:29]),
		.chany_top_in(sb_1__1__33_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__32_ccff_tail),
		.chany_bottom_out(cby_1__1__37_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__37_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__37_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__37_ccff_tail));

	cby_1__1_ cby_5__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__33_chany_top_out[0:29]),
		.chany_top_in(sb_1__1__34_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__33_ccff_tail),
		.chany_bottom_out(cby_1__1__38_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__38_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__38_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__38_ccff_tail));

	cby_1__1_ cby_5__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__34_chany_top_out[0:29]),
		.chany_top_in(sb_1__8__4_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__34_ccff_tail),
		.chany_bottom_out(cby_1__1__39_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__39_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__39_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__39_ccff_tail));

	cby_1__1_ cby_6__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__0__5_chany_top_out[0:29]),
		.chany_top_in(sb_1__1__35_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__0__5_ccff_tail),
		.chany_bottom_out(cby_1__1__40_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__40_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__40_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__40_ccff_tail));

	cby_1__1_ cby_6__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__35_chany_top_out[0:29]),
		.chany_top_in(sb_1__1__36_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__35_ccff_tail),
		.chany_bottom_out(cby_1__1__41_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__41_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__41_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__41_ccff_tail));

	cby_1__1_ cby_6__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__36_chany_top_out[0:29]),
		.chany_top_in(sb_1__1__37_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__36_ccff_tail),
		.chany_bottom_out(cby_1__1__42_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__42_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__42_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__42_ccff_tail));

	cby_1__1_ cby_6__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__37_chany_top_out[0:29]),
		.chany_top_in(sb_1__1__38_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__37_ccff_tail),
		.chany_bottom_out(cby_1__1__43_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__43_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__43_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__43_ccff_tail));

	cby_1__1_ cby_6__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__38_chany_top_out[0:29]),
		.chany_top_in(sb_1__1__39_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__38_ccff_tail),
		.chany_bottom_out(cby_1__1__44_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__44_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__44_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__44_ccff_tail));

	cby_1__1_ cby_6__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__39_chany_top_out[0:29]),
		.chany_top_in(sb_1__1__40_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__39_ccff_tail),
		.chany_bottom_out(cby_1__1__45_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__45_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__45_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__45_ccff_tail));

	cby_1__1_ cby_6__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__40_chany_top_out[0:29]),
		.chany_top_in(sb_1__1__41_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__40_ccff_tail),
		.chany_bottom_out(cby_1__1__46_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__46_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__46_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__46_ccff_tail));

	cby_1__1_ cby_6__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__41_chany_top_out[0:29]),
		.chany_top_in(sb_1__8__5_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__41_ccff_tail),
		.chany_bottom_out(cby_1__1__47_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__47_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__47_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__47_ccff_tail));

	cby_1__1_ cby_7__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__0__6_chany_top_out[0:29]),
		.chany_top_in(sb_1__1__42_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__0__6_ccff_tail),
		.chany_bottom_out(cby_1__1__48_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__48_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__48_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__48_ccff_tail));

	cby_1__1_ cby_7__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__42_chany_top_out[0:29]),
		.chany_top_in(sb_1__1__43_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__42_ccff_tail),
		.chany_bottom_out(cby_1__1__49_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__49_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__49_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__49_ccff_tail));

	cby_1__1_ cby_7__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__43_chany_top_out[0:29]),
		.chany_top_in(sb_1__1__44_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__43_ccff_tail),
		.chany_bottom_out(cby_1__1__50_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__50_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__50_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__50_ccff_tail));

	cby_1__1_ cby_7__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__44_chany_top_out[0:29]),
		.chany_top_in(sb_1__1__45_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__44_ccff_tail),
		.chany_bottom_out(cby_1__1__51_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__51_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__51_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__51_ccff_tail));

	cby_1__1_ cby_7__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__45_chany_top_out[0:29]),
		.chany_top_in(sb_1__1__46_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__45_ccff_tail),
		.chany_bottom_out(cby_1__1__52_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__52_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__52_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__52_ccff_tail));

	cby_1__1_ cby_7__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__46_chany_top_out[0:29]),
		.chany_top_in(sb_1__1__47_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__46_ccff_tail),
		.chany_bottom_out(cby_1__1__53_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__53_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__53_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__53_ccff_tail));

	cby_1__1_ cby_7__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__47_chany_top_out[0:29]),
		.chany_top_in(sb_1__1__48_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__47_ccff_tail),
		.chany_bottom_out(cby_1__1__54_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__54_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__54_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__54_ccff_tail));

	cby_1__1_ cby_7__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_1__1__48_chany_top_out[0:29]),
		.chany_top_in(sb_1__8__6_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__48_ccff_tail),
		.chany_bottom_out(cby_1__1__55_chany_bottom_out[0:29]),
		.chany_top_out(cby_1__1__55_chany_top_out[0:29]),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_1__1__55_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_1__1__55_ccff_tail));

	cby_8__1_ cby_8__1_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_8__0__0_chany_top_out[0:29]),
		.chany_top_in(sb_8__1__0_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__0__7_ccff_tail),
		.chany_bottom_out(cby_8__1__0_chany_bottom_out[0:29]),
		.chany_top_out(cby_8__1__0_chany_top_out[0:29]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_8__1__0_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_8__1__0_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_8__1__0_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_8__1__0_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_8__1__0_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_8__1__0_ccff_tail));

	cby_8__1_ cby_8__2_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_8__1__0_chany_top_out[0:29]),
		.chany_top_in(sb_8__1__1_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__49_ccff_tail),
		.chany_bottom_out(cby_8__1__1_chany_bottom_out[0:29]),
		.chany_top_out(cby_8__1__1_chany_top_out[0:29]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_8__1__1_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_8__1__1_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_8__1__1_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_8__1__1_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_8__1__1_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_8__1__1_ccff_tail));

	cby_8__1_ cby_8__3_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_8__1__1_chany_top_out[0:29]),
		.chany_top_in(sb_8__1__2_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__50_ccff_tail),
		.chany_bottom_out(cby_8__1__2_chany_bottom_out[0:29]),
		.chany_top_out(cby_8__1__2_chany_top_out[0:29]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_8__1__2_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_8__1__2_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_8__1__2_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_8__1__2_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_8__1__2_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_8__1__2_ccff_tail));

	cby_8__1_ cby_8__4_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_8__1__2_chany_top_out[0:29]),
		.chany_top_in(sb_8__1__3_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__51_ccff_tail),
		.chany_bottom_out(cby_8__1__3_chany_bottom_out[0:29]),
		.chany_top_out(cby_8__1__3_chany_top_out[0:29]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_8__1__3_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_8__1__3_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_8__1__3_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_8__1__3_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_8__1__3_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_8__1__3_ccff_tail));

	cby_8__1_ cby_8__5_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_8__1__3_chany_top_out[0:29]),
		.chany_top_in(sb_8__1__4_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__52_ccff_tail),
		.chany_bottom_out(cby_8__1__4_chany_bottom_out[0:29]),
		.chany_top_out(cby_8__1__4_chany_top_out[0:29]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_8__1__4_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_8__1__4_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_8__1__4_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_8__1__4_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_8__1__4_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_8__1__4_ccff_tail));

	cby_8__1_ cby_8__6_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_8__1__4_chany_top_out[0:29]),
		.chany_top_in(sb_8__1__5_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__53_ccff_tail),
		.chany_bottom_out(cby_8__1__5_chany_bottom_out[0:29]),
		.chany_top_out(cby_8__1__5_chany_top_out[0:29]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_8__1__5_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_8__1__5_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_8__1__5_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_8__1__5_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_8__1__5_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_8__1__5_ccff_tail));

	cby_8__1_ cby_8__7_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_8__1__5_chany_top_out[0:29]),
		.chany_top_in(sb_8__1__6_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__54_ccff_tail),
		.chany_bottom_out(cby_8__1__6_chany_bottom_out[0:29]),
		.chany_top_out(cby_8__1__6_chany_top_out[0:29]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_8__1__6_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_8__1__6_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_8__1__6_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_8__1__6_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_8__1__6_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_8__1__6_ccff_tail));

	cby_8__1_ cby_8__8_ (
		.pReset(pReset),
		.prog_clk(prog_clk),
		.chany_bottom_in(sb_8__1__6_chany_top_out[0:29]),
		.chany_top_in(sb_8__8__0_chany_bottom_out[0:29]),
		.ccff_head(cbx_1__1__55_ccff_tail),
		.chany_bottom_out(cby_8__1__7_chany_bottom_out[0:29]),
		.chany_top_out(cby_8__1__7_chany_top_out[0:29]),
		.right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_(cby_8__1__7_right_grid_left_width_0_height_0_subtile_0__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_(cby_8__1__7_right_grid_left_width_0_height_0_subtile_1__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_(cby_8__1__7_right_grid_left_width_0_height_0_subtile_2__pin_outpad_0_),
		.right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_(cby_8__1__7_right_grid_left_width_0_height_0_subtile_3__pin_outpad_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_0_(cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I4_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4_1_(cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I4_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_(cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I4i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_(cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I4i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_0_(cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I5_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5_1_(cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I5_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_(cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I5i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_(cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I5i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_0_(cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I6_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6_1_(cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I6_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_(cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I6i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_(cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I6i_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_0_(cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I7_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7_1_(cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I7_1_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_(cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I7i_0_),
		.left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_(cby_8__1__7_left_grid_right_width_0_height_0_subtile_0__pin_I7i_1_),
		.ccff_tail(cby_8__1__7_ccff_tail));

	direct_interc direct_interc_0_ (
		.in(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_0_out));

	direct_interc direct_interc_1_ (
		.in(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_1_out));

	direct_interc direct_interc_2_ (
		.in(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_2_out));

	direct_interc direct_interc_3_ (
		.in(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_3_out));

	direct_interc direct_interc_4_ (
		.in(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_4_out));

	direct_interc direct_interc_5_ (
		.in(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_5_out));

	direct_interc direct_interc_6_ (
		.in(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_6_out));

	direct_interc direct_interc_7_ (
		.in(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_7_out));

	direct_interc direct_interc_8_ (
		.in(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_8_out));

	direct_interc direct_interc_9_ (
		.in(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_9_out));

	direct_interc direct_interc_10_ (
		.in(grid_clb_12_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_10_out));

	direct_interc direct_interc_11_ (
		.in(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_11_out));

	direct_interc direct_interc_12_ (
		.in(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_12_out));

	direct_interc direct_interc_13_ (
		.in(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_13_out));

	direct_interc direct_interc_14_ (
		.in(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_14_out));

	direct_interc direct_interc_15_ (
		.in(grid_clb_18_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_15_out));

	direct_interc direct_interc_16_ (
		.in(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_16_out));

	direct_interc direct_interc_17_ (
		.in(grid_clb_20_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_17_out));

	direct_interc direct_interc_18_ (
		.in(grid_clb_21_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_18_out));

	direct_interc direct_interc_19_ (
		.in(grid_clb_22_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_19_out));

	direct_interc direct_interc_20_ (
		.in(grid_clb_23_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_20_out));

	direct_interc direct_interc_21_ (
		.in(grid_clb_25_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_21_out));

	direct_interc direct_interc_22_ (
		.in(grid_clb_26_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_22_out));

	direct_interc direct_interc_23_ (
		.in(grid_clb_27_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_23_out));

	direct_interc direct_interc_24_ (
		.in(grid_clb_28_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_24_out));

	direct_interc direct_interc_25_ (
		.in(grid_clb_29_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_25_out));

	direct_interc direct_interc_26_ (
		.in(grid_clb_30_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_26_out));

	direct_interc direct_interc_27_ (
		.in(grid_clb_31_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_27_out));

	direct_interc direct_interc_28_ (
		.in(grid_clb_33_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_28_out));

	direct_interc direct_interc_29_ (
		.in(grid_clb_34_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_29_out));

	direct_interc direct_interc_30_ (
		.in(grid_clb_35_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_30_out));

	direct_interc direct_interc_31_ (
		.in(grid_clb_36_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_31_out));

	direct_interc direct_interc_32_ (
		.in(grid_clb_37_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_32_out));

	direct_interc direct_interc_33_ (
		.in(grid_clb_38_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_33_out));

	direct_interc direct_interc_34_ (
		.in(grid_clb_39_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_34_out));

	direct_interc direct_interc_35_ (
		.in(grid_clb_41_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_35_out));

	direct_interc direct_interc_36_ (
		.in(grid_clb_42_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_36_out));

	direct_interc direct_interc_37_ (
		.in(grid_clb_43_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_37_out));

	direct_interc direct_interc_38_ (
		.in(grid_clb_44_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_38_out));

	direct_interc direct_interc_39_ (
		.in(grid_clb_45_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_39_out));

	direct_interc direct_interc_40_ (
		.in(grid_clb_46_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_40_out));

	direct_interc direct_interc_41_ (
		.in(grid_clb_47_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_41_out));

	direct_interc direct_interc_42_ (
		.in(grid_clb_49_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_42_out));

	direct_interc direct_interc_43_ (
		.in(grid_clb_50_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_43_out));

	direct_interc direct_interc_44_ (
		.in(grid_clb_51_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_44_out));

	direct_interc direct_interc_45_ (
		.in(grid_clb_52_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_45_out));

	direct_interc direct_interc_46_ (
		.in(grid_clb_53_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_46_out));

	direct_interc direct_interc_47_ (
		.in(grid_clb_54_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_47_out));

	direct_interc direct_interc_48_ (
		.in(grid_clb_55_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_48_out));

	direct_interc direct_interc_49_ (
		.in(grid_clb_57_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_49_out));

	direct_interc direct_interc_50_ (
		.in(grid_clb_58_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_50_out));

	direct_interc direct_interc_51_ (
		.in(grid_clb_59_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_51_out));

	direct_interc direct_interc_52_ (
		.in(grid_clb_60_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_52_out));

	direct_interc direct_interc_53_ (
		.in(grid_clb_61_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_53_out));

	direct_interc direct_interc_54_ (
		.in(grid_clb_62_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_54_out));

	direct_interc direct_interc_55_ (
		.in(grid_clb_63_bottom_width_0_height_0_subtile_0__pin_cout_0_),
		.out(direct_interc_55_out));

	direct_interc direct_interc_56_ (
		.in(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_56_out));

	direct_interc direct_interc_57_ (
		.in(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_57_out));

	direct_interc direct_interc_58_ (
		.in(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_58_out));

	direct_interc direct_interc_59_ (
		.in(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_59_out));

	direct_interc direct_interc_60_ (
		.in(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_60_out));

	direct_interc direct_interc_61_ (
		.in(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_61_out));

	direct_interc direct_interc_62_ (
		.in(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_62_out));

	direct_interc direct_interc_63_ (
		.in(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_63_out));

	direct_interc direct_interc_64_ (
		.in(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_64_out));

	direct_interc direct_interc_65_ (
		.in(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_65_out));

	direct_interc direct_interc_66_ (
		.in(grid_clb_12_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_66_out));

	direct_interc direct_interc_67_ (
		.in(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_67_out));

	direct_interc direct_interc_68_ (
		.in(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_68_out));

	direct_interc direct_interc_69_ (
		.in(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_69_out));

	direct_interc direct_interc_70_ (
		.in(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_70_out));

	direct_interc direct_interc_71_ (
		.in(grid_clb_18_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_71_out));

	direct_interc direct_interc_72_ (
		.in(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_72_out));

	direct_interc direct_interc_73_ (
		.in(grid_clb_20_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_73_out));

	direct_interc direct_interc_74_ (
		.in(grid_clb_21_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_74_out));

	direct_interc direct_interc_75_ (
		.in(grid_clb_22_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_75_out));

	direct_interc direct_interc_76_ (
		.in(grid_clb_23_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_76_out));

	direct_interc direct_interc_77_ (
		.in(grid_clb_25_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_77_out));

	direct_interc direct_interc_78_ (
		.in(grid_clb_26_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_78_out));

	direct_interc direct_interc_79_ (
		.in(grid_clb_27_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_79_out));

	direct_interc direct_interc_80_ (
		.in(grid_clb_28_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_80_out));

	direct_interc direct_interc_81_ (
		.in(grid_clb_29_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_81_out));

	direct_interc direct_interc_82_ (
		.in(grid_clb_30_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_82_out));

	direct_interc direct_interc_83_ (
		.in(grid_clb_31_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_83_out));

	direct_interc direct_interc_84_ (
		.in(grid_clb_33_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_84_out));

	direct_interc direct_interc_85_ (
		.in(grid_clb_34_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_85_out));

	direct_interc direct_interc_86_ (
		.in(grid_clb_35_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_86_out));

	direct_interc direct_interc_87_ (
		.in(grid_clb_36_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_87_out));

	direct_interc direct_interc_88_ (
		.in(grid_clb_37_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_88_out));

	direct_interc direct_interc_89_ (
		.in(grid_clb_38_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_89_out));

	direct_interc direct_interc_90_ (
		.in(grid_clb_39_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_90_out));

	direct_interc direct_interc_91_ (
		.in(grid_clb_41_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_91_out));

	direct_interc direct_interc_92_ (
		.in(grid_clb_42_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_92_out));

	direct_interc direct_interc_93_ (
		.in(grid_clb_43_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_93_out));

	direct_interc direct_interc_94_ (
		.in(grid_clb_44_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_94_out));

	direct_interc direct_interc_95_ (
		.in(grid_clb_45_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_95_out));

	direct_interc direct_interc_96_ (
		.in(grid_clb_46_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_96_out));

	direct_interc direct_interc_97_ (
		.in(grid_clb_47_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_97_out));

	direct_interc direct_interc_98_ (
		.in(grid_clb_49_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_98_out));

	direct_interc direct_interc_99_ (
		.in(grid_clb_50_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_99_out));

	direct_interc direct_interc_100_ (
		.in(grid_clb_51_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_100_out));

	direct_interc direct_interc_101_ (
		.in(grid_clb_52_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_101_out));

	direct_interc direct_interc_102_ (
		.in(grid_clb_53_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_102_out));

	direct_interc direct_interc_103_ (
		.in(grid_clb_54_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_103_out));

	direct_interc direct_interc_104_ (
		.in(grid_clb_55_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_104_out));

	direct_interc direct_interc_105_ (
		.in(grid_clb_57_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_105_out));

	direct_interc direct_interc_106_ (
		.in(grid_clb_58_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_106_out));

	direct_interc direct_interc_107_ (
		.in(grid_clb_59_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_107_out));

	direct_interc direct_interc_108_ (
		.in(grid_clb_60_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_108_out));

	direct_interc direct_interc_109_ (
		.in(grid_clb_61_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_109_out));

	direct_interc direct_interc_110_ (
		.in(grid_clb_62_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_110_out));

	direct_interc direct_interc_111_ (
		.in(grid_clb_63_bottom_width_0_height_0_subtile_0__pin_reg_out_0_),
		.out(direct_interc_111_out));

	direct_interc direct_interc_112_ (
		.in(grid_clb_1_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_112_out));

	direct_interc direct_interc_113_ (
		.in(grid_clb_2_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_113_out));

	direct_interc direct_interc_114_ (
		.in(grid_clb_3_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_114_out));

	direct_interc direct_interc_115_ (
		.in(grid_clb_4_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_115_out));

	direct_interc direct_interc_116_ (
		.in(grid_clb_5_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_116_out));

	direct_interc direct_interc_117_ (
		.in(grid_clb_6_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_117_out));

	direct_interc direct_interc_118_ (
		.in(grid_clb_7_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_118_out));

	direct_interc direct_interc_119_ (
		.in(grid_clb_9_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_119_out));

	direct_interc direct_interc_120_ (
		.in(grid_clb_10_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_120_out));

	direct_interc direct_interc_121_ (
		.in(grid_clb_11_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_121_out));

	direct_interc direct_interc_122_ (
		.in(grid_clb_12_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_122_out));

	direct_interc direct_interc_123_ (
		.in(grid_clb_13_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_123_out));

	direct_interc direct_interc_124_ (
		.in(grid_clb_14_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_124_out));

	direct_interc direct_interc_125_ (
		.in(grid_clb_15_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_125_out));

	direct_interc direct_interc_126_ (
		.in(grid_clb_17_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_126_out));

	direct_interc direct_interc_127_ (
		.in(grid_clb_18_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_127_out));

	direct_interc direct_interc_128_ (
		.in(grid_clb_19_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_128_out));

	direct_interc direct_interc_129_ (
		.in(grid_clb_20_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_129_out));

	direct_interc direct_interc_130_ (
		.in(grid_clb_21_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_130_out));

	direct_interc direct_interc_131_ (
		.in(grid_clb_22_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_131_out));

	direct_interc direct_interc_132_ (
		.in(grid_clb_23_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_132_out));

	direct_interc direct_interc_133_ (
		.in(grid_clb_25_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_133_out));

	direct_interc direct_interc_134_ (
		.in(grid_clb_26_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_134_out));

	direct_interc direct_interc_135_ (
		.in(grid_clb_27_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_135_out));

	direct_interc direct_interc_136_ (
		.in(grid_clb_28_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_136_out));

	direct_interc direct_interc_137_ (
		.in(grid_clb_29_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_137_out));

	direct_interc direct_interc_138_ (
		.in(grid_clb_30_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_138_out));

	direct_interc direct_interc_139_ (
		.in(grid_clb_31_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_139_out));

	direct_interc direct_interc_140_ (
		.in(grid_clb_33_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_140_out));

	direct_interc direct_interc_141_ (
		.in(grid_clb_34_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_141_out));

	direct_interc direct_interc_142_ (
		.in(grid_clb_35_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_142_out));

	direct_interc direct_interc_143_ (
		.in(grid_clb_36_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_143_out));

	direct_interc direct_interc_144_ (
		.in(grid_clb_37_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_144_out));

	direct_interc direct_interc_145_ (
		.in(grid_clb_38_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_145_out));

	direct_interc direct_interc_146_ (
		.in(grid_clb_39_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_146_out));

	direct_interc direct_interc_147_ (
		.in(grid_clb_41_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_147_out));

	direct_interc direct_interc_148_ (
		.in(grid_clb_42_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_148_out));

	direct_interc direct_interc_149_ (
		.in(grid_clb_43_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_149_out));

	direct_interc direct_interc_150_ (
		.in(grid_clb_44_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_150_out));

	direct_interc direct_interc_151_ (
		.in(grid_clb_45_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_151_out));

	direct_interc direct_interc_152_ (
		.in(grid_clb_46_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_152_out));

	direct_interc direct_interc_153_ (
		.in(grid_clb_47_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_153_out));

	direct_interc direct_interc_154_ (
		.in(grid_clb_49_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_154_out));

	direct_interc direct_interc_155_ (
		.in(grid_clb_50_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_155_out));

	direct_interc direct_interc_156_ (
		.in(grid_clb_51_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_156_out));

	direct_interc direct_interc_157_ (
		.in(grid_clb_52_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_157_out));

	direct_interc direct_interc_158_ (
		.in(grid_clb_53_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_158_out));

	direct_interc direct_interc_159_ (
		.in(grid_clb_54_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_159_out));

	direct_interc direct_interc_160_ (
		.in(grid_clb_55_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_160_out));

	direct_interc direct_interc_161_ (
		.in(grid_clb_57_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_161_out));

	direct_interc direct_interc_162_ (
		.in(grid_clb_58_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_162_out));

	direct_interc direct_interc_163_ (
		.in(grid_clb_59_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_163_out));

	direct_interc direct_interc_164_ (
		.in(grid_clb_60_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_164_out));

	direct_interc direct_interc_165_ (
		.in(grid_clb_61_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_165_out));

	direct_interc direct_interc_166_ (
		.in(grid_clb_62_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_166_out));

	direct_interc direct_interc_167_ (
		.in(grid_clb_63_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_167_out));

	direct_interc direct_interc_168_ (
		.in(grid_clb_0_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_168_out));

	direct_interc direct_interc_169_ (
		.in(grid_clb_8_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_169_out));

	direct_interc direct_interc_170_ (
		.in(grid_clb_16_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_170_out));

	direct_interc direct_interc_171_ (
		.in(grid_clb_24_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_171_out));

	direct_interc direct_interc_172_ (
		.in(grid_clb_32_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_172_out));

	direct_interc direct_interc_173_ (
		.in(grid_clb_40_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_173_out));

	direct_interc direct_interc_174_ (
		.in(grid_clb_48_bottom_width_0_height_0_subtile_0__pin_sc_out_0_),
		.out(direct_interc_174_out));

endmodule
// ----- END Verilog module for fpga_top -----

//----- Default net type -----
`default_nettype none




