//-------------------------------------------
//	FPGA Synthesizable Verilog Netlist
//	Description: Verilog netlist for pre-configured FPGA fabric by design: maskmul
//	Author: Xifan TANG
//	Organization: University of Utah
//	Date: Thu Dec  5 17:13:01 2024
//-------------------------------------------
//----- Time scale -----
`timescale 1ns / 1ps

//----- Default net type -----
`default_nettype wire

module maskmul_top_formal_verification (
input [0:0] am_0_,
input [0:0] am_1_,
input [0:0] bm_0_,
input [0:0] bm_1_,
input [0:0] ma_0_,
input [0:0] ma_1_,
input [0:0] mb_0_,
input [0:0] mb_1_,
input [0:0] mq_0_,
input [0:0] mq_1_,
input [0:0] reset,
input [0:0] clock,
output [0:0] qm_0_,
output [0:0] qm_1_);

// ----- Local wires for FPGA fabric -----
wire [0:0] clk_fm;
wire [0:0] reset_fm;
wire [0:127] gfpga_pad_io_soc_in_fm;
wire [0:127] gfpga_pad_io_soc_out_fm;
wire [0:127] gfpga_pad_io_soc_dir_fm;
wire [0:0] ccff_head_fm;
wire [0:0] ccff_tail_fm;
wire [0:0] isol_n_fm;
wire [0:0] prog_reset_fm;
wire [0:0] prog_clk_fm;
wire [0:0] test_enable_fm;

// ----- FPGA top-level module to be capsulated -----
	fpga_top U0_formal_verification (
		clk_fm[0],
		reset_fm[0],
		isol_n_fm[0],
		prog_reset_fm[0],
		prog_clk_fm[0],
		test_enable_fm[0],
		gfpga_pad_io_soc_in_fm[0:127],
		gfpga_pad_io_soc_out_fm[0:127],
		gfpga_pad_io_soc_dir_fm[0:127],
		ccff_head_fm[0],
		ccff_tail_fm[0]);

// ----- Begin Connect Global ports of FPGA top module -----
	assign test_enable_fm[0] = 1'b0;
	assign prog_clk_fm[0] = 1'b0;
	assign prog_reset_fm[0] = 1'b1;
	assign isol_n_fm[0] = 1'b1;
	assign clk_fm[0] = clock[0];
	assign reset_fm[0] = 1'b1;
// ----- End Connect Global ports of FPGA top module -----

// ----- Link BLIF Benchmark I/Os to FPGA I/Os -----
// ----- Blif Benchmark input am_0_ is mapped to FPGA IOPAD gfpga_pad_io_soc_in_fm[49] -----
	assign gfpga_pad_io_soc_in_fm[49] = am_0_[0];

// ----- Blif Benchmark input am_1_ is mapped to FPGA IOPAD gfpga_pad_io_soc_in_fm[48] -----
	assign gfpga_pad_io_soc_in_fm[48] = am_1_[0];

// ----- Blif Benchmark input bm_0_ is mapped to FPGA IOPAD gfpga_pad_io_soc_in_fm[51] -----
	assign gfpga_pad_io_soc_in_fm[51] = bm_0_[0];

// ----- Blif Benchmark input bm_1_ is mapped to FPGA IOPAD gfpga_pad_io_soc_in_fm[50] -----
	assign gfpga_pad_io_soc_in_fm[50] = bm_1_[0];

// ----- Blif Benchmark input ma_0_ is mapped to FPGA IOPAD gfpga_pad_io_soc_in_fm[53] -----
	assign gfpga_pad_io_soc_in_fm[53] = ma_0_[0];

// ----- Blif Benchmark input ma_1_ is mapped to FPGA IOPAD gfpga_pad_io_soc_in_fm[52] -----
	assign gfpga_pad_io_soc_in_fm[52] = ma_1_[0];

// ----- Blif Benchmark input mb_0_ is mapped to FPGA IOPAD gfpga_pad_io_soc_in_fm[55] -----
	assign gfpga_pad_io_soc_in_fm[55] = mb_0_[0];

// ----- Blif Benchmark input mb_1_ is mapped to FPGA IOPAD gfpga_pad_io_soc_in_fm[54] -----
	assign gfpga_pad_io_soc_in_fm[54] = mb_1_[0];

// ----- Blif Benchmark input mq_0_ is mapped to FPGA IOPAD gfpga_pad_io_soc_in_fm[57] -----
	assign gfpga_pad_io_soc_in_fm[57] = mq_0_[0];

// ----- Blif Benchmark input mq_1_ is mapped to FPGA IOPAD gfpga_pad_io_soc_in_fm[56] -----
	assign gfpga_pad_io_soc_in_fm[56] = mq_1_[0];

// ----- Blif Benchmark input reset is mapped to FPGA IOPAD gfpga_pad_io_soc_in_fm[60] -----
	assign gfpga_pad_io_soc_in_fm[60] = reset[0];

// ----- Blif Benchmark input clock is mapped to FPGA IOPAD gfpga_pad_io_soc_in_fm[61] -----
	assign gfpga_pad_io_soc_in_fm[61] = clock[0];

// ----- Blif Benchmark output qm_0_ is mapped to FPGA IOPAD gfpga_pad_io_soc_out_fm[59] -----
	assign qm_0_[0] = gfpga_pad_io_soc_out_fm[59];

// ----- Blif Benchmark output qm_1_ is mapped to FPGA IOPAD gfpga_pad_io_soc_out_fm[58] -----
	assign qm_1_[0] = gfpga_pad_io_soc_out_fm[58];

// ----- Wire unused FPGA I/Os to constants -----
	assign gfpga_pad_io_soc_in_fm[0] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[1] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[2] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[3] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[4] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[5] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[6] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[7] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[8] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[9] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[10] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[11] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[12] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[13] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[14] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[15] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[16] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[17] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[18] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[19] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[20] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[21] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[22] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[23] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[24] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[25] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[26] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[27] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[28] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[29] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[30] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[31] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[32] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[33] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[34] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[35] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[36] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[37] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[38] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[39] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[40] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[41] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[42] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[43] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[44] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[45] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[46] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[47] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[58] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[59] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[62] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[63] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[64] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[65] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[66] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[67] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[68] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[69] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[70] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[71] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[72] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[73] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[74] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[75] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[76] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[77] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[78] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[79] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[80] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[81] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[82] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[83] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[84] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[85] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[86] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[87] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[88] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[89] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[90] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[91] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[92] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[93] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[94] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[95] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[96] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[97] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[98] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[99] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[100] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[101] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[102] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[103] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[104] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[105] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[106] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[107] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[108] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[109] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[110] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[111] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[112] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[113] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[114] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[115] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[116] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[117] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[118] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[119] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[120] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[121] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[122] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[123] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[124] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[125] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[126] = 1'b0;
	assign gfpga_pad_io_soc_in_fm[127] = 1'b0;


// ----- Begin load bitstream to configuration memories -----
// ----- Begin assign bitstream to configuration memories -----
initial begin
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_1__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_2__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_3__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_4__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_5__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_6__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_7__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__1_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__2_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = 17'b00111100000000001;
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = 2'b01;
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = 2'b01;
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = 2'b01;
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = 17'b00010010000000001;
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = 2'b01;
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = 2'b01;
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = 17'b00111100000000001;
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = 2'b01;
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = 2'b01;
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = 2'b01;
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = 17'b10100110011010100;
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = 2'b01;
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = 2'b01;
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = 17'b00000110011000000;
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = 2'b01;
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = 2'b01;
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = 17'b00010100001010000;
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = 2'b01;
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = 2'b01;
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = 17'b00010010010010000;
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = 2'b01;
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = 2'b01;
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = 17'b00001001000001100;
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = 2'b01;
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.grid_clb_8__3_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__4_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__5_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__6_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__7_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_1.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_2.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_3.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_4.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_5.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_6.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_mode_default__frac_lut4_0.frac_lut4_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0:16] = {17{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_logic_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.logical_tile_clb_mode_default__fle_mode_physical__fabric_mode_default__frac_logic_0.mem_frac_lut4_0_in_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_fabric_out_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_0_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_clb_8__8_.logical_tile_clb_mode_clb__0.logical_tile_clb_mode_default__fle_7.logical_tile_clb_mode_default__fle_mode_physical__fabric_0.mem_ff_1_D_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.grid_io_top_top_1__9_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_top_1__9_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_top_1__9_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_top_1__9_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_top_2__9_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_top_2__9_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_top_2__9_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_top_2__9_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_top_3__9_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_top_3__9_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_top_3__9_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_top_3__9_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_top_4__9_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_top_4__9_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_top_4__9_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_top_4__9_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_top_5__9_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_top_5__9_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_top_5__9_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_top_5__9_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_top_6__9_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_top_6__9_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_top_6__9_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_top_6__9_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_top_7__9_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_top_7__9_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_top_7__9_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_top_7__9_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_top_8__9_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_top_8__9_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_top_8__9_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_top_top_8__9_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_right_9__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_right_9__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_right_9__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_right_9__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_right_9__7_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_right_9__7_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_right_9__7_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_right_9__7_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_right_9__6_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_right_9__6_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_right_9__6_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_right_9__6_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_right_9__5_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_right_9__5_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_right_9__5_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_right_9__5_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_right_9__4_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_right_9__4_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_right_9__4_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_right_9__4_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_right_9__3_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_right_9__3_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_right_9__3_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_right_9__3_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_right_9__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_right_9__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_right_9__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_right_9__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b0;
	force U0_formal_verification.grid_io_right_right_9__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_right_9__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_right_9__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_right_right_9__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_bottom_8__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_bottom_7__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_bottom_7__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_bottom_7__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_bottom_7__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_bottom_6__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_bottom_6__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_bottom_6__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_bottom_6__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_bottom_5__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_bottom_5__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_bottom_5__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_bottom_5__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_bottom_4__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_bottom_4__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_bottom_4__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_bottom_4__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_bottom_3__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_bottom_3__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_bottom_3__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_bottom_3__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_bottom_2__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_bottom_2__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_bottom_2__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_bottom_2__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_bottom_1__0_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_bottom_1__0_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_bottom_1__0_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_bottom_bottom_1__0_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_left_0__1_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_left_0__1_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_left_0__1_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_left_0__1_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_left_0__2_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_left_0__2_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_left_0__2_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_left_0__2_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_left_0__3_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_left_0__3_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_left_0__3_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_left_0__3_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_left_0__4_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_left_0__4_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_left_0__4_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_left_0__4_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_left_0__5_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_left_0__5_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_left_0__5_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_left_0__5_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_left_0__6_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_left_0__6_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_left_0__6_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_left_0__6_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_left_0__7_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_left_0__7_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_left_0__7_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_left_0__7_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_left_0__8_.logical_tile_io_mode_io__0.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_left_0__8_.logical_tile_io_mode_io__1.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_left_0__8_.logical_tile_io_mode_io__2.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.grid_io_left_left_0__8_.logical_tile_io_mode_io__3.logical_tile_io_mode_physical__iopad_0.io_sky130_fd_sc_hd__dfrtp_1_mem.mem_out[0] = 1'b1;
	force U0_formal_verification.sb_0__0_.mem_top_track_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_4.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_6.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_8.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_10.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_12.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_14.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_16.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_18.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_28.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_46.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_48.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_top_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_0.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_2.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_4.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_6.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_8.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_10.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_12.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_14.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_16.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_18.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_28.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_46.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_48.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__0_.mem_right_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_top_track_2.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_top_track_4.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_top_track_6.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_top_track_10.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_top_track_12.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_top_track_20.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_top_track_28.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_top_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_2.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_4.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_6.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_10.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_12.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_14.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_18.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_20.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_22.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_24.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_26.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_28.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_38.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_40.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_46.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_48.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_52.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_54.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_right_track_56.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_3.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_5.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_7.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_11.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_13.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_21.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_29.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__1_.mem_bottom_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_2.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_4.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_6.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_10.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_12.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_20.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_28.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_2.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_4.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_6.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_10.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_12.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_14.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_18.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_20.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_22.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_24.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_26.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_28.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_38.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_40.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_46.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_48.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_52.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_54.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_right_track_56.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_3.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_5.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_7.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_11.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_13.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_21.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_29.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__2_.mem_bottom_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_2.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_4.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_6.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_10.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_12.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_20.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_28.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_2.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_4.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_6.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_10.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_12.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_14.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_18.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_20.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_22.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_24.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_26.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_28.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_38.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_40.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_46.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_48.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_52.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_54.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_right_track_56.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_3.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_5.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_7.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_11.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_13.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_21.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_29.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__3_.mem_bottom_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_2.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_4.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_6.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_10.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_12.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_20.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_28.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_2.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_4.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_6.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_10.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_12.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_14.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_18.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_20.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_22.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_24.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_26.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_28.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_38.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_40.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_46.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_48.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_52.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_54.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_right_track_56.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_3.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_5.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_7.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_11.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_13.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_21.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_29.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__4_.mem_bottom_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_2.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_4.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_6.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_10.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_12.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_20.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_28.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_2.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_4.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_6.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_10.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_12.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_14.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_18.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_20.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_22.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_24.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_26.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_28.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_38.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_40.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_46.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_48.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_52.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_54.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_right_track_56.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_3.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_5.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_7.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_11.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_13.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_21.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_29.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__5_.mem_bottom_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_top_track_2.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_top_track_4.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_top_track_6.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_top_track_10.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_top_track_12.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_top_track_20.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_top_track_28.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_top_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_2.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_4.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_6.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_10.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_12.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_14.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_18.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_20.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_22.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_24.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_26.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_28.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_38.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_40.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_46.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_48.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_52.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_54.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_right_track_56.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_3.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_5.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_7.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_11.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_13.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_21.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_29.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__6_.mem_bottom_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_top_track_2.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_top_track_4.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_top_track_6.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_top_track_10.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_top_track_12.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_top_track_20.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_top_track_28.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_top_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_2.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_4.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_6.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_10.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_12.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_14.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_18.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_20.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_22.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_24.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_26.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_28.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_38.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_40.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_46.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_48.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_52.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_54.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_right_track_56.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_3.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_5.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_7.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_11.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_13.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_21.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_29.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__7_.mem_bottom_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_2.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_4.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_6.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_10.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_12.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_14.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_16.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_18.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_20.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_22.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_24.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_26.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_28.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_36.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_38.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_40.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_42.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_46.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_48.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_52.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_54.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_56.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_right_track_58.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_17.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_19.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_0__8_.mem_bottom_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_2.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_4.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_6.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_10.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_12.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_14.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_18.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_20.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_22.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_24.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_26.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_28.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_36.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_40.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_42.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_46.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_48.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_top_track_58.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_2.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_4.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_6.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_10.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_12.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_20.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_28.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_right_track_52.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_3.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_5.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_7.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_11.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_13.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_21.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_29.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__0_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_top_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_top_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_top_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_top_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__1_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__2_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__3_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__4_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__5_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_top_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_top_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_top_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_top_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__6_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_top_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_top_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_top_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_top_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_right_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_right_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__7_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_right_track_12.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_right_track_20.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_right_track_28.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_3.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_5.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_7.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_11.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_13.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_15.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_19.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_21.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_bottom_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_left_track_13.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_left_track_21.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_left_track_29.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_1__8_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_2.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_4.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_6.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_10.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_12.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_14.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_18.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_20.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_22.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_24.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_26.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_28.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_36.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_40.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_42.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_46.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_48.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_top_track_58.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_2.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_4.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_6.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_10.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_12.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_20.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_28.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_right_track_52.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_3.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_5.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_7.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_11.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_13.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_21.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_29.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__0_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__1_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_right_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_right_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__2_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__3_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__4_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__5_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_top_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_top_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_top_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_top_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__6_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_top_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_top_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_top_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_top_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_right_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_right_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__7_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_right_track_12.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_right_track_20.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_right_track_28.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_3.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_5.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_7.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_11.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_13.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_15.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_19.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_21.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_bottom_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_left_track_13.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_left_track_21.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_left_track_29.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_2__8_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_2.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_4.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_6.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_10.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_12.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_14.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_18.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_20.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_22.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_24.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_26.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_28.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_36.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_40.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_42.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_46.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_48.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_top_track_58.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_2.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_4.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_6.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_10.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_12.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_20.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_28.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_right_track_52.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_3.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_5.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_7.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_11.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_13.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_21.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_29.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__0_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_top_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_top_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_top_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_top_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__1_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__2_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__3_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__4_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__5_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_top_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_top_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_top_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_top_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__6_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_top_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_top_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_top_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_top_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_right_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_right_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__7_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_right_track_12.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_right_track_20.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_right_track_28.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_3.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_5.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_7.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_11.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_13.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_15.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_19.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_21.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_bottom_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_left_track_13.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_left_track_21.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_left_track_29.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_3__8_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_2.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_4.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_6.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_10.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_12.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_14.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_18.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_20.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_22.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_24.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_26.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_28.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_36.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_40.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_42.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_46.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_48.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_top_track_58.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_right_track_2.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_right_track_4.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_right_track_6.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_right_track_10.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_right_track_12.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_right_track_20.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_right_track_28.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_right_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_right_track_52.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_3.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_5.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_7.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_11.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_13.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_21.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_29.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__0_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_right_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_right_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__1_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_right_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_right_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__2_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_right_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_right_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__3_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_right_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_right_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__4_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_right_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_right_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__5_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_top_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_top_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_top_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_top_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_right_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_right_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__6_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_top_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_top_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_top_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_top_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_right_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_right_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__7_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_right_track_12.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_right_track_20.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_right_track_28.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_3.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_5.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_7.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_11.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_13.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_15.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_19.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_21.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_bottom_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_left_track_13.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_left_track_21.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_left_track_29.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_4__8_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_2.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_4.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_6.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_10.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_12.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_14.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_18.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_20.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_22.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_24.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_26.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_28.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_36.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_5__0_.mem_top_track_40.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_42.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_46.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_48.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_top_track_58.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_right_track_2.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_right_track_4.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_right_track_6.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_right_track_10.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_right_track_12.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_right_track_20.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_right_track_28.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_right_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_right_track_52.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_left_track_3.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_left_track_5.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_left_track_7.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_left_track_11.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_left_track_13.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_left_track_21.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_left_track_29.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__0_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_top_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_top_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_top_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_top_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_right_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_right_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__1_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_top_track_0.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_5__2_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_top_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_top_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_top_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_top_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_right_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_right_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__2_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_top_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_top_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_top_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_top_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_right_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_right_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_right_track_44.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_5__3_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__3_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_top_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_top_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_top_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_top_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_right_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_right_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__4_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_top_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_top_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_top_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_top_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_right_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_right_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__5_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_top_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_top_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_top_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_top_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_right_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_right_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_bottom_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_bottom_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_bottom_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__6_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_top_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_top_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_top_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_top_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_right_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_right_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__7_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_right_track_12.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_right_track_20.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_right_track_28.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_3.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_5.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_7.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_11.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_13.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_15.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_19.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_21.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_bottom_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_left_track_13.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_left_track_21.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_left_track_29.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_5__8_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_2.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_4.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_6.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_10.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_12.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_14.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_18.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_20.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_22.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_24.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_26.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_28.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_36.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_40.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_42.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_46.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_48.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_top_track_58.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_right_track_2.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_right_track_4.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_right_track_6.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_right_track_10.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_right_track_12.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_right_track_20.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_right_track_28.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_right_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_right_track_52.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_left_track_3.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_left_track_5.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_left_track_7.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_left_track_11.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_left_track_13.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_left_track_21.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_left_track_29.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__0_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_top_track_4.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__1_.mem_top_track_6.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_6__1_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_top_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_top_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_top_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_right_track_12.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_6__1_.mem_right_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_right_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__1_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_top_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_top_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_top_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_top_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_right_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_right_track_28.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_6__2_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__2_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_top_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_top_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_top_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_top_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_right_track_20.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_6__3_.mem_right_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_21.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_6__3_.mem_bottom_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__3_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_top_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_top_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_top_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_top_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_right_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_right_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__4_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_top_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_top_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_top_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_top_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_right_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_right_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__5_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_top_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_top_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_top_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_top_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_right_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_right_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_bottom_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_bottom_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_bottom_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__6_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_top_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_top_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_top_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_top_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_right_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_right_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__7_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_right_track_12.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_right_track_20.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_right_track_28.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_3.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_5.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_7.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_11.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_13.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_15.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_19.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_21.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_bottom_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_left_track_13.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_left_track_21.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_left_track_29.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_6__8_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_2.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_4.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_6.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_10.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_12.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_7__0_.mem_top_track_14.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_16.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_18.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_20.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_22.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_24.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_26.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_28.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_36.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_40.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_42.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_44.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_46.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_48.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_top_track_58.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_right_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_right_track_2.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_right_track_4.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_right_track_6.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_right_track_10.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_right_track_12.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_right_track_20.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_7__0_.mem_right_track_28.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_right_track_44.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_7__0_.mem_right_track_52.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_3.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_5.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_7.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_11.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_13.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_21.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_29.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__0_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_top_track_6.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_7__1_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_top_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_top_track_20.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_7__1_.mem_top_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_top_track_44.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_7__1_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_right_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_right_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__1_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_top_track_4.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_7__2_.mem_top_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_top_track_12.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_7__2_.mem_top_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_top_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_right_track_2.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_7__2_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_right_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_right_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__2_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_top_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_top_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_top_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_top_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_right_track_0.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_7__3_.mem_right_track_2.mem_out[0:3] = 4'b1001;
	force U0_formal_verification.sb_7__3_.mem_right_track_4.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.sb_7__3_.mem_right_track_6.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_7__3_.mem_right_track_10.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_7__3_.mem_right_track_12.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_7__3_.mem_right_track_20.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_7__3_.mem_right_track_28.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_7__3_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_13.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_7__3_.mem_bottom_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_29.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_7__3_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__3_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_top_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_top_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_top_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_top_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_right_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_right_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__4_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_top_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_top_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_top_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_top_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_right_track_0.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_7__5_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_right_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_right_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_37.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_7__5_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__5_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_top_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_top_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_top_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_top_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_right_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_right_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__6_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_top_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_top_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_top_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_top_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_right_track_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_right_track_20.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_right_track_28.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_21.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_29.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__7_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_right_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_right_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_right_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_right_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_right_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_right_track_12.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_right_track_20.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_right_track_28.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_right_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_right_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_right_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_3.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_5.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_7.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_11.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_13.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_15.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_19.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_21.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_bottom_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_left_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_left_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_left_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_left_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_left_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_left_track_13.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_left_track_21.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_left_track_29.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_left_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_left_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_7__8_.mem_left_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_0.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_2.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_4.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_6.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_8.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_10.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_12.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_14.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_16.mem_out[0:1] = 2'b10;
	force U0_formal_verification.sb_8__0_.mem_top_track_18.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_20.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_22.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_24.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_26.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_28.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_top_track_30.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_32.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_34.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_36.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_38.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_40.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_8__0_.mem_top_track_42.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_44.mem_out[0:1] = 2'b01;
	force U0_formal_verification.sb_8__0_.mem_top_track_46.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_48.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_top_track_50.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_left_track_1.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_left_track_3.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_left_track_5.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_left_track_7.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_left_track_9.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_left_track_11.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_left_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_left_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_left_track_17.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_left_track_19.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_left_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_left_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_left_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_left_track_35.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__0_.mem_left_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_left_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_left_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__0_.mem_left_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_top_track_6.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_8__1_.mem_top_track_10.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_8__1_.mem_top_track_12.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_top_track_20.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_top_track_28.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_13.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_21.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_29.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_left_track_3.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_left_track_5.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_left_track_7.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_left_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_left_track_11.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_left_track_13.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_left_track_15.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_8__1_.mem_left_track_17.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_left_track_19.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_left_track_21.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_left_track_23.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_left_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_left_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_left_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_left_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_left_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_left_track_35.mem_out[0:1] = {2{1'b1}};
	force U0_formal_verification.sb_8__1_.mem_left_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_left_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_left_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_left_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_left_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_left_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_left_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_left_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__1_.mem_left_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_top_track_2.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_8__2_.mem_top_track_4.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.sb_8__2_.mem_top_track_6.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_8__2_.mem_top_track_10.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.sb_8__2_.mem_top_track_12.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_top_track_20.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_top_track_28.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_8__2_.mem_top_track_36.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_8__2_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_top_track_52.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_8__2_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_bottom_track_3.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_8__2_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_bottom_track_7.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.sb_8__2_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_bottom_track_13.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_bottom_track_21.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_bottom_track_29.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_left_track_3.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_left_track_5.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_left_track_7.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_left_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_left_track_11.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_left_track_13.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_left_track_15.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_left_track_19.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_left_track_21.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_left_track_23.mem_out[0:2] = {3{1'b1}};
	force U0_formal_verification.sb_8__2_.mem_left_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_left_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_left_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_left_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_left_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_left_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_left_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_left_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_left_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_left_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_left_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_left_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_left_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_left_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__2_.mem_left_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_top_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_top_track_12.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_top_track_20.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_top_track_28.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_bottom_track_1.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_8__3_.mem_bottom_track_3.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_8__3_.mem_bottom_track_5.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_8__3_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_bottom_track_11.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.sb_8__3_.mem_bottom_track_13.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_8__3_.mem_bottom_track_21.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_8__3_.mem_bottom_track_29.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_8__3_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_bottom_track_53.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_8__3_.mem_left_track_1.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_8__3_.mem_left_track_3.mem_out[0:2] = 3'b010;
	force U0_formal_verification.sb_8__3_.mem_left_track_5.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_8__3_.mem_left_track_7.mem_out[0:2] = 3'b110;
	force U0_formal_verification.sb_8__3_.mem_left_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_left_track_11.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_8__3_.mem_left_track_13.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_left_track_15.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_left_track_19.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_left_track_21.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_left_track_23.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_left_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_left_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_left_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_left_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_left_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_left_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_left_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_left_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_left_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_left_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_left_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_left_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_left_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_left_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__3_.mem_left_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_top_track_0.mem_out[0:3] = 4'b0001;
	force U0_formal_verification.sb_8__4_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_top_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_top_track_12.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_top_track_20.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_top_track_28.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_7.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.sb_8__4_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_13.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_8__4_.mem_bottom_track_21.mem_out[0:2] = 3'b101;
	force U0_formal_verification.sb_8__4_.mem_bottom_track_29.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_37.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_8__4_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_left_track_3.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_left_track_5.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_left_track_7.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_left_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_left_track_11.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_left_track_13.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_left_track_15.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_left_track_19.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_left_track_21.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_left_track_23.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_left_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_left_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_left_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_left_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_left_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_left_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_left_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_left_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_left_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_left_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_left_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_left_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_left_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_left_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__4_.mem_left_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_top_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_top_track_12.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_top_track_20.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_top_track_28.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_13.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_21.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_29.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_bottom_track_53.mem_out[0:2] = 3'b001;
	force U0_formal_verification.sb_8__5_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_left_track_3.mem_out[0:2] = 3'b011;
	force U0_formal_verification.sb_8__5_.mem_left_track_5.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_left_track_7.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_left_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_left_track_11.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_left_track_13.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_left_track_15.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_left_track_19.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_left_track_21.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_left_track_23.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_left_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_left_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_left_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_left_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_left_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_left_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_left_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_left_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_left_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_left_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_left_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_left_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_left_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_left_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__5_.mem_left_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_top_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_top_track_12.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_top_track_20.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_top_track_28.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_bottom_track_13.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_bottom_track_21.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_bottom_track_29.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_left_track_3.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_left_track_5.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_left_track_7.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_left_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_left_track_11.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_left_track_13.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_left_track_15.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_left_track_19.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_left_track_21.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_left_track_23.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_left_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_left_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_left_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_left_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_left_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_left_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_left_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_left_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_left_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_left_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_left_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_left_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_left_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_left_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__6_.mem_left_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_top_track_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_top_track_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_top_track_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_top_track_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_top_track_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_top_track_12.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_top_track_20.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_top_track_28.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_top_track_36.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_top_track_44.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_top_track_52.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_13.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_21.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_29.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_37.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_45.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_bottom_track_53.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_3.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_5.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_7.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_11.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_13.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_15.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_17.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_19.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_21.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_23.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__7_.mem_left_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_3.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_5.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_7.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_11.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_17.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_19.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_21.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_bottom_track_59.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_1.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_3.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_5.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_7.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_9.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_11.mem_out[0:2] = {3{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_13.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_15.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_17.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_19.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_21.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_23.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_25.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_27.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_29.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_31.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_33.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_35.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_37.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_39.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_41.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_43.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_45.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_47.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_49.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_51.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_53.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_55.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_57.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.sb_8__8_.mem_left_track_59.mem_out[0:1] = {2{1'b0}};
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__0_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__1_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__2_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__3_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__3_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__3_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__3_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__3_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__3_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__3_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__3_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__3_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__3_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__3_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__3_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__3_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__3_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__3_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__3_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__4_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__5_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__6_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__6_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__6_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__6_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__6_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__6_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__6_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__6_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__6_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__6_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__6_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__6_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__6_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__6_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__6_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__6_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__7_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__7_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__7_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__7_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__7_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__7_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__7_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__7_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__7_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__7_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__7_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__7_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__7_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__7_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__7_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__7_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__8_.mem_bottom_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__8_.mem_bottom_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__8_.mem_bottom_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__8_.mem_bottom_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__8_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__8_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__8_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__8_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__8_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__8_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__8_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__8_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__8_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__8_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__8_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__8_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__8_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__8_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__8_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_1__8_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__0_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__1_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__1_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__1_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__1_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__1_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__1_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__1_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__1_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__1_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__1_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__1_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__1_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__1_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__1_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__1_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__1_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__2_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__3_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__3_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__3_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__3_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__3_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__3_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__3_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__3_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__3_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__3_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__3_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__3_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__3_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__3_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__3_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__3_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__4_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__4_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__4_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__4_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__4_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__4_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__4_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__4_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__4_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__4_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__4_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__4_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__4_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__4_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__4_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__4_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__5_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__5_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__5_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__5_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__5_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__5_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__5_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__5_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__5_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__5_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__5_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__5_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__5_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__5_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__5_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__5_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__6_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__6_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__6_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__6_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__6_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__6_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__6_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__6_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__6_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__6_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__6_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__6_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__6_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__6_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__6_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__6_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__7_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__7_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__7_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__7_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__7_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__7_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__7_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__7_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__7_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__7_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__7_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__7_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__7_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__7_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__7_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__7_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__8_.mem_bottom_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__8_.mem_bottom_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__8_.mem_bottom_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__8_.mem_bottom_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__8_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__8_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__8_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__8_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__8_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__8_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__8_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__8_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__8_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__8_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__8_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__8_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__8_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__8_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__8_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_2__8_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__0_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__1_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__1_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__1_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__1_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__1_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__1_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__1_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__1_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__1_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__1_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__1_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__1_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__1_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__1_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__1_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__1_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__2_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__3_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__3_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__3_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__3_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__3_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__3_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__3_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__3_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__3_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__3_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__3_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__3_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__3_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__3_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__3_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__3_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__4_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__4_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__4_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__4_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__4_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__4_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__4_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__4_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__4_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__4_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__4_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__4_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__4_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__4_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__4_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__4_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__5_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__5_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__5_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__5_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__5_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__5_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__5_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__5_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__5_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__5_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__5_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__5_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__5_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__5_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__5_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__5_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__6_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__6_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__6_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__6_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__6_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__6_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__6_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__6_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__6_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__6_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__6_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__6_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__6_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__6_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__6_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__6_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__7_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__7_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__7_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__7_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__7_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__7_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__7_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__7_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__7_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__7_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__7_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__7_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__7_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__7_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__7_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__7_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__8_.mem_bottom_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__8_.mem_bottom_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__8_.mem_bottom_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__8_.mem_bottom_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__8_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__8_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__8_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__8_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__8_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__8_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__8_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__8_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__8_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__8_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__8_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__8_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__8_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__8_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__8_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_3__8_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__0_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__1_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__2_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__3_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__3_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__3_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__3_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__3_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__3_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__3_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__3_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__3_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__3_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__3_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__3_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__3_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__3_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__3_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__3_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__4_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__5_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__6_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__6_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__6_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__6_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__6_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__6_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__6_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__6_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__6_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__6_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__6_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__6_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__6_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__6_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__6_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__6_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__7_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__7_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__7_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__7_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__7_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__7_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__7_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__7_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__7_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__7_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__7_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__7_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__7_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__7_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__7_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__7_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__8_.mem_bottom_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__8_.mem_bottom_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__8_.mem_bottom_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__8_.mem_bottom_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__8_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__8_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__8_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__8_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__8_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__8_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__8_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__8_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__8_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__8_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__8_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__8_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__8_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__8_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__8_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_4__8_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__0_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__0_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__0_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__0_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__1_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__2_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__2_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__2_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__2_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__2_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__2_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__2_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__2_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__2_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__2_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__2_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__2_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__2_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__2_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__2_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__2_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__3_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__3_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__3_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__3_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__3_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__3_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__3_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__3_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__3_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__3_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__3_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__3_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__3_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__3_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__3_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__3_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__4_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__4_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__4_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__4_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__4_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__4_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__4_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__4_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__4_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__4_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__4_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__4_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__4_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__4_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__4_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__4_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__5_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__5_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__5_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__5_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__5_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__5_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__5_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__5_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__5_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__5_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__5_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__5_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__5_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__5_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__5_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__5_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__6_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__6_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__6_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__6_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__6_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__6_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__6_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__6_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__6_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__6_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__6_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__6_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__6_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__6_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__6_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__6_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__7_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__7_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__7_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__7_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__7_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__7_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__7_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__7_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__7_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__7_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__7_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__7_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__7_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__7_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__7_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__7_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__8_.mem_bottom_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__8_.mem_bottom_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__8_.mem_bottom_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__8_.mem_bottom_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__8_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__8_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__8_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__8_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__8_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__8_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__8_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__8_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__8_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__8_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__8_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__8_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__8_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__8_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__8_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_5__8_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__0_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__0_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__0_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__0_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__1_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__1_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__1_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__1_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__1_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__1_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__1_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__1_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__1_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__1_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__1_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__1_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__1_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__1_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__1_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__1_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__2_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__2_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__2_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__2_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__2_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__2_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__2_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__2_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__2_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__2_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__2_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__2_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__2_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__2_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__2_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__2_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__3_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__3_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__3_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__3_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__3_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__3_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__3_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__3_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__3_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__3_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__3_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__3_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__3_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__3_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__3_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__3_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__4_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__4_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__4_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__4_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__4_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__4_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__4_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__4_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__4_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__4_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__4_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__4_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__4_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__4_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__4_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__4_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__5_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__5_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__5_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__5_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__5_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__5_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__5_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__5_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__5_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__5_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__5_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__5_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__5_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__5_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__5_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__5_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__6_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__7_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__7_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__7_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__7_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__7_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__7_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__7_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__7_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__7_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__7_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__7_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__7_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__7_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__7_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__7_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__7_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__8_.mem_bottom_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__8_.mem_bottom_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__8_.mem_bottom_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__8_.mem_bottom_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__8_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__8_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__8_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__8_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__8_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__8_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__8_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__8_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__8_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__8_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__8_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__8_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__8_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__8_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__8_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_6__8_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__0_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__0_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__0_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__0_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__1_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__1_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__1_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__1_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__1_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__1_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__1_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__1_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__1_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__1_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__1_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__1_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__1_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__1_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__1_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__1_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__2_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__2_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__2_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__2_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__2_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__2_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__2_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__2_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__2_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__2_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__2_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__2_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__2_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__2_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__2_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__2_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__3_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__3_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__3_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__3_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__3_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__3_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__3_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__3_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__3_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__3_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__3_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__3_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__3_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__3_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__3_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__3_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__4_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__4_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__4_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__4_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__4_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__4_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__4_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__4_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__4_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__4_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__4_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__4_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__4_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__4_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__4_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__4_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__5_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__5_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__5_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__5_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__5_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__5_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__5_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__5_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__5_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__5_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__5_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__5_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__5_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__5_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__5_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__5_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__6_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__6_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__6_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__6_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__6_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__6_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__6_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__6_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__6_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__6_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__6_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__6_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__6_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__6_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__6_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__6_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__7_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__7_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__7_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__7_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__7_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__7_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__7_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__7_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__7_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__7_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__7_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__7_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__7_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__7_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__7_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__7_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__8_.mem_bottom_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__8_.mem_bottom_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__8_.mem_bottom_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__8_.mem_bottom_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__8_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__8_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__8_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__8_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__8_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__8_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__8_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__8_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__8_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__8_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__8_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__8_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__8_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__8_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__8_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_7__8_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__0_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__0_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__0_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__0_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__1_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__1_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__1_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__1_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__1_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__1_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__1_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__1_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__1_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__1_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__1_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__1_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__1_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__1_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__1_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__1_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__2_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__2_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__2_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__2_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__2_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__2_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__2_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__2_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__2_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__2_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__2_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__2_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__2_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__2_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__2_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__2_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__3_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__3_.mem_top_ipin_1.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_8__3_.mem_top_ipin_2.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.cbx_8__3_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__3_.mem_top_ipin_4.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.cbx_8__3_.mem_top_ipin_5.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.cbx_8__3_.mem_top_ipin_6.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.cbx_8__3_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__3_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__3_.mem_top_ipin_9.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.cbx_8__3_.mem_top_ipin_10.mem_out[0:3] = 4'b1101;
	force U0_formal_verification.cbx_8__3_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__3_.mem_top_ipin_12.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.cbx_8__3_.mem_top_ipin_13.mem_out[0:3] = 4'b0110;
	force U0_formal_verification.cbx_8__3_.mem_top_ipin_14.mem_out[0:3] = 4'b1001;
	force U0_formal_verification.cbx_8__3_.mem_top_ipin_15.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.cbx_8__4_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__4_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__4_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__4_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__4_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__4_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__4_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__4_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__4_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__4_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__4_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__4_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__4_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__4_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__4_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__4_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__5_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__5_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__5_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__5_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__5_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__5_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__5_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__5_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__5_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__5_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__5_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__5_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__5_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__5_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__5_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__5_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__6_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__6_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__6_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__6_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__6_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__6_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__6_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__6_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__6_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__6_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__6_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__6_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__6_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__6_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__6_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__6_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__7_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__7_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__7_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__7_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__7_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__7_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__7_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__7_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__7_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__7_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__7_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__7_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__7_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__7_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__7_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__7_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__8_.mem_bottom_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__8_.mem_bottom_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__8_.mem_bottom_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__8_.mem_bottom_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__8_.mem_top_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__8_.mem_top_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__8_.mem_top_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__8_.mem_top_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__8_.mem_top_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__8_.mem_top_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__8_.mem_top_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__8_.mem_top_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__8_.mem_top_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__8_.mem_top_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__8_.mem_top_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__8_.mem_top_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__8_.mem_top_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__8_.mem_top_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__8_.mem_top_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cbx_8__8_.mem_top_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_0__1_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_0__1_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_0__1_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_0__1_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_0__2_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_0__3_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_0__3_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_0__3_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_0__3_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_0__4_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_0__4_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_0__4_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_0__4_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_0__5_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_0__6_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_0__6_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_0__6_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_0__6_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_0__7_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_0__7_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_0__7_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_0__7_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_0__8_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_0__8_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_0__8_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_0__8_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__1_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__2_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__3_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__3_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__3_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__3_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__3_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__3_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__3_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__3_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__3_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__3_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__3_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__3_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__3_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__3_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__3_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__3_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__4_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__4_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__4_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__4_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__4_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__4_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__4_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__4_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__4_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__4_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__4_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__4_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__4_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__4_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__4_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__4_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__5_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__6_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__6_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__6_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__6_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__6_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__6_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__6_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__6_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__6_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__6_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__6_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__6_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__6_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__6_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__6_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__6_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__7_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__7_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__7_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__7_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__7_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__7_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__7_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__7_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__7_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__7_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__7_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__7_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__7_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__7_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__7_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__7_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__8_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__8_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__8_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__8_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__8_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__8_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__8_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__8_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__8_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__8_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__8_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__8_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__8_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__8_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__8_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_1__8_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__1_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__2_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__2_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__2_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__2_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__2_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__2_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__2_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__2_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__2_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__2_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__2_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__2_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__2_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__2_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__2_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__2_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__3_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__3_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__3_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__3_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__3_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__3_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__3_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__3_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__3_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__3_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__3_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__3_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__3_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__3_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__3_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__3_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__4_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__4_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__4_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__4_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__4_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__4_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__4_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__4_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__4_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__4_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__4_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__4_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__4_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__4_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__4_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__4_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__5_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__5_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__5_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__5_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__5_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__5_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__5_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__5_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__5_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__5_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__5_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__5_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__5_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__5_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__5_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__5_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__6_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__6_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__6_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__6_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__6_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__6_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__6_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__6_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__6_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__6_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__6_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__6_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__6_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__6_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__6_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__6_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__7_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__7_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__7_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__7_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__7_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__7_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__7_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__7_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__7_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__7_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__7_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__7_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__7_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__7_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__7_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__7_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__8_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__8_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__8_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__8_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__8_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__8_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__8_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__8_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__8_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__8_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__8_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__8_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__8_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__8_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__8_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_2__8_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__1_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__1_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__1_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__1_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__1_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__1_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__1_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__1_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__1_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__1_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__1_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__1_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__1_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__1_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__1_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__1_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__2_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__3_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__3_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__3_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__3_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__3_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__3_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__3_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__3_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__3_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__3_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__3_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__3_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__3_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__3_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__3_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__3_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__4_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__4_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__4_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__4_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__4_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__4_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__4_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__4_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__4_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__4_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__4_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__4_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__4_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__4_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__4_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__4_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__5_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__6_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__6_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__6_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__6_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__6_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__6_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__6_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__6_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__6_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__6_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__6_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__6_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__6_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__6_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__6_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__6_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__7_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__7_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__7_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__7_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__7_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__7_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__7_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__7_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__7_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__7_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__7_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__7_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__7_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__7_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__7_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__7_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__8_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__8_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__8_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__8_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__8_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__8_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__8_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__8_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__8_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__8_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__8_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__8_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__8_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__8_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__8_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_3__8_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__1_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__1_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__1_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__1_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__1_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__1_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__1_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__1_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__1_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__1_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__1_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__1_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__1_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__1_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__1_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__1_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__2_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__3_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__3_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__3_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__3_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__3_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__3_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__3_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__3_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__3_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__3_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__3_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__3_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__3_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__3_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__3_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__3_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__4_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__4_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__4_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__4_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__4_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__4_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__4_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__4_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__4_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__4_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__4_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__4_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__4_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__4_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__4_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__4_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__5_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__6_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__6_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__6_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__6_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__6_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__6_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__6_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__6_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__6_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__6_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__6_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__6_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__6_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__6_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__6_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__6_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__7_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__7_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__7_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__7_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__7_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__7_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__7_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__7_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__7_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__7_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__7_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__7_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__7_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__7_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__7_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__7_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__8_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__8_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__8_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__8_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__8_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__8_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__8_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__8_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__8_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__8_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__8_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__8_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__8_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__8_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__8_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_4__8_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__1_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__1_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__1_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__1_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__1_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__1_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__1_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__1_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__1_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__1_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__1_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__1_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__1_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__1_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__1_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__1_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__2_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__2_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__2_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__2_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__2_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__2_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__2_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__2_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__2_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__2_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__2_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__2_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__2_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__2_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__2_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__2_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__3_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__3_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__3_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__3_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__3_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__3_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__3_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__3_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__3_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__3_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__3_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__3_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__3_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__3_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__3_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__3_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__4_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__4_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__4_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__4_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__4_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__4_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__4_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__4_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__4_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__4_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__4_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__4_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__4_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__4_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__4_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__4_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__5_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__5_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__5_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__5_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__5_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__5_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__5_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__5_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__5_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__5_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__5_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__5_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__5_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__5_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__5_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__5_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__6_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__6_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__6_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__6_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__6_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__6_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__6_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__6_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__6_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__6_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__6_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__6_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__6_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__6_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__6_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__6_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__7_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__7_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__7_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__7_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__7_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__7_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__7_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__7_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__7_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__7_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__7_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__7_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__7_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__7_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__7_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__7_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__8_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__8_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__8_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__8_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__8_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__8_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__8_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__8_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__8_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__8_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__8_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__8_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__8_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__8_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__8_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_5__8_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__1_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__1_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__1_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__1_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__1_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__1_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__1_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__1_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__1_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__1_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__1_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__1_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__1_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__1_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__1_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__1_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__2_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__2_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__2_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__2_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__2_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__2_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__2_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__2_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__2_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__2_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__2_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__2_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__2_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__2_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__2_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__2_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__3_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__3_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__3_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__3_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__3_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__3_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__3_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__3_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__3_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__3_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__3_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__3_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__3_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__3_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__3_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__3_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__4_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__4_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__4_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__4_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__4_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__4_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__4_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__4_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__4_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__4_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__4_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__4_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__4_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__4_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__4_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__4_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__5_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__5_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__5_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__5_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__5_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__5_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__5_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__5_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__5_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__5_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__5_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__5_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__5_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__5_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__5_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__5_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__6_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__6_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__6_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__6_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__6_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__6_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__6_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__6_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__6_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__6_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__6_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__6_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__6_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__6_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__6_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__6_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__7_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__7_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__7_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__7_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__7_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__7_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__7_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__7_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__7_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__7_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__7_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__7_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__7_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__7_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__7_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__7_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__8_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__8_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__8_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__8_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__8_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__8_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__8_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__8_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__8_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__8_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__8_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__8_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__8_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__8_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__8_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_6__8_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__1_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__1_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__1_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__1_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__1_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__1_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__1_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__1_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__1_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__1_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__1_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__1_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__1_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__1_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__1_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__1_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__2_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__2_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__2_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__2_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__2_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__2_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__2_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__2_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__2_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__2_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__2_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__2_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__2_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__2_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__2_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__2_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__3_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__3_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__3_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__3_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__3_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__3_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__3_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__3_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__3_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__3_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__3_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__3_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__3_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__3_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__3_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__3_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__4_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__4_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__4_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__4_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__4_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__4_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__4_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__4_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__4_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__4_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__4_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__4_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__4_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__4_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__4_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__4_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__5_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__5_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__5_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__5_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__5_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__5_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__5_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__5_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__5_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__5_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__5_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__5_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__5_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__5_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__5_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__5_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__6_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__6_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__6_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__6_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__6_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__6_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__6_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__6_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__6_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__6_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__6_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__6_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__6_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__6_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__6_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__6_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__7_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__7_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__7_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__7_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__7_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__7_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__7_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__7_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__7_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__7_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__7_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__7_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__7_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__7_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__7_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__7_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__8_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__8_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__8_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__8_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__8_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__8_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__8_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__8_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__8_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__8_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__8_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__8_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__8_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__8_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__8_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_7__8_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__1_.mem_left_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__1_.mem_left_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__1_.mem_left_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__1_.mem_left_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__1_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__1_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__1_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__1_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__1_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__1_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__1_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__1_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__1_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__1_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__1_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__1_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__1_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__1_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__1_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__1_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__2_.mem_left_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__2_.mem_left_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__2_.mem_left_ipin_2.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.cby_8__2_.mem_left_ipin_3.mem_out[0:3] = 4'b1110;
	force U0_formal_verification.cby_8__2_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__2_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__2_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__2_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__2_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__2_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__2_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__2_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__2_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__2_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__2_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__2_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__2_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__2_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__2_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__2_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__3_.mem_left_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__3_.mem_left_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__3_.mem_left_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__3_.mem_left_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__3_.mem_right_ipin_0.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.cby_8__3_.mem_right_ipin_1.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.cby_8__3_.mem_right_ipin_2.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.cby_8__3_.mem_right_ipin_3.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.cby_8__3_.mem_right_ipin_4.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.cby_8__3_.mem_right_ipin_5.mem_out[0:3] = 4'b0111;
	force U0_formal_verification.cby_8__3_.mem_right_ipin_6.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.cby_8__3_.mem_right_ipin_7.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.cby_8__3_.mem_right_ipin_8.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.cby_8__3_.mem_right_ipin_9.mem_out[0:3] = 4'b0011;
	force U0_formal_verification.cby_8__3_.mem_right_ipin_10.mem_out[0:3] = 4'b1001;
	force U0_formal_verification.cby_8__3_.mem_right_ipin_11.mem_out[0:3] = 4'b1011;
	force U0_formal_verification.cby_8__3_.mem_right_ipin_12.mem_out[0:3] = 4'b0100;
	force U0_formal_verification.cby_8__3_.mem_right_ipin_13.mem_out[0:3] = {4{1'b1}};
	force U0_formal_verification.cby_8__3_.mem_right_ipin_14.mem_out[0:3] = 4'b0010;
	force U0_formal_verification.cby_8__3_.mem_right_ipin_15.mem_out[0:3] = 4'b0101;
	force U0_formal_verification.cby_8__4_.mem_left_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__4_.mem_left_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__4_.mem_left_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__4_.mem_left_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__4_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__4_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__4_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__4_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__4_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__4_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__4_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__4_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__4_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__4_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__4_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__4_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__4_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__4_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__4_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__4_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__5_.mem_left_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__5_.mem_left_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__5_.mem_left_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__5_.mem_left_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__5_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__5_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__5_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__5_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__5_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__5_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__5_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__5_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__5_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__5_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__5_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__5_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__5_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__5_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__5_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__5_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__6_.mem_left_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__6_.mem_left_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__6_.mem_left_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__6_.mem_left_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__6_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__6_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__6_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__6_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__6_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__6_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__6_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__6_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__6_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__6_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__6_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__6_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__6_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__6_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__6_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__6_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__7_.mem_left_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__7_.mem_left_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__7_.mem_left_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__7_.mem_left_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__7_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__7_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__7_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__7_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__7_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__7_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__7_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__7_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__7_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__7_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__7_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__7_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__7_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__7_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__7_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__7_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__8_.mem_left_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__8_.mem_left_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__8_.mem_left_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__8_.mem_left_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__8_.mem_right_ipin_0.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__8_.mem_right_ipin_1.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__8_.mem_right_ipin_2.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__8_.mem_right_ipin_3.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__8_.mem_right_ipin_4.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__8_.mem_right_ipin_5.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__8_.mem_right_ipin_6.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__8_.mem_right_ipin_7.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__8_.mem_right_ipin_8.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__8_.mem_right_ipin_9.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__8_.mem_right_ipin_10.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__8_.mem_right_ipin_11.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__8_.mem_right_ipin_12.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__8_.mem_right_ipin_13.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__8_.mem_right_ipin_14.mem_out[0:3] = {4{1'b0}};
	force U0_formal_verification.cby_8__8_.mem_right_ipin_15.mem_out[0:3] = {4{1'b0}};
end
// ----- End assign bitstream to configuration memories -----
// ----- End load bitstream to configuration memories -----
endmodule
// ----- END Verilog module for maskmul_top_formal_verification -----

//----- Default net type -----
`default_nettype none

